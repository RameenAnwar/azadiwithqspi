##
## LEF for PtnCells ;
## created by Innovus v20.10-p004_1 on Sat May 28 13:30:04 2022
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO azadi_soc_top_caravel
  CLASS BLOCK ;
  SIZE 2399.820000 BY 2599.980000 ;
  FOREIGN azadi_soc_top_caravel 0.000000 0.000000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 319.264 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 1596.09 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 4.795000 0.000000 4.935000 0.490000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 41.5651 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 207.546 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAPARTIALMETALAREA 0.255 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.808 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 6.1578 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 33.312 LAYER met4  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.495 LAYER met4  ;
    ANTENNAMAXAREACAR 68.182 LAYER met4  ;
    ANTENNAMAXSIDEAREACAR 345.881 LAYER met4  ;
    ANTENNAMAXCUTCAR 0.265455 LAYER via4  ;
    PORT
      LAYER met2 ;
        RECT 0.000000 1.120000 0.485000 1.260000 ;
    END
  END wb_rst_i
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.100000 0.000000 506.240000 0.490000 ;
    END
  END wbs_stb_i
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.275000 0.000000 170.415000 0.490000 ;
    END
  END wbs_cyc_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 510.965000 0.000000 511.105000 0.490000 ;
    END
  END wbs_we_i
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.230000 0.000000 501.370000 0.490000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.365000 0.000000 496.505000 0.490000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.495000 0.000000 491.635000 0.490000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.630000 0.000000 486.770000 0.490000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.020000 0.000000 326.160000 0.490000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.150000 0.000000 321.290000 0.490000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.285000 0.000000 316.425000 0.490000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 311.420000 0.000000 311.560000 0.490000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.550000 0.000000 306.690000 0.490000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.685000 0.000000 301.825000 0.490000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.815000 0.000000 296.955000 0.490000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.950000 0.000000 292.090000 0.490000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.085000 0.000000 287.225000 0.490000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 282.215000 0.000000 282.355000 0.490000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.350000 0.000000 277.490000 0.490000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.480000 0.000000 272.620000 0.490000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.615000 0.000000 267.755000 0.490000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750000 0.000000 262.890000 0.490000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.880000 0.000000 258.020000 0.490000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.015000 0.000000 253.155000 0.490000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.145000 0.000000 248.285000 0.490000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.280000 0.000000 243.420000 0.490000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.415000 0.000000 238.555000 0.490000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.545000 0.000000 233.685000 0.490000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.680000 0.000000 228.820000 0.490000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.810000 0.000000 223.950000 0.490000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.945000 0.000000 219.085000 0.490000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.080000 0.000000 214.220000 0.490000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.210000 0.000000 209.350000 0.490000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.345000 0.000000 204.485000 0.490000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.475000 0.000000 199.615000 0.490000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.610000 0.000000 194.750000 0.490000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.745000 0.000000 189.885000 0.490000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.875000 0.000000 185.015000 0.490000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.010000 0.000000 180.150000 0.490000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.140000 0.000000 175.280000 0.490000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.410000 0.000000 165.550000 0.490000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.540000 0.000000 160.680000 0.490000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.675000 0.000000 155.815000 0.490000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.805000 0.000000 150.945000 0.490000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.940000 0.000000 146.080000 0.490000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.075000 0.000000 141.215000 0.490000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.205000 0.000000 136.345000 0.490000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.340000 0.000000 131.480000 0.490000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.470000 0.000000 126.610000 0.490000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.605000 0.000000 121.745000 0.490000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.740000 0.000000 116.880000 0.490000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 111.870000 0.000000 112.010000 0.490000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.005000 0.000000 107.145000 0.490000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.135000 0.000000 102.275000 0.490000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.270000 0.000000 97.410000 0.490000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.405000 0.000000 92.545000 0.490000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.535000 0.000000 87.675000 0.490000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.670000 0.000000 82.810000 0.490000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.800000 0.000000 77.940000 0.490000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 72.935000 0.000000 73.075000 0.490000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.070000 0.000000 68.210000 0.490000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.200000 0.000000 63.340000 0.490000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.335000 0.000000 58.475000 0.490000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.465000 0.000000 53.605000 0.490000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.600000 0.000000 48.740000 0.490000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.735000 0.000000 43.875000 0.490000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.865000 0.000000 39.005000 0.490000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.000000 0.000000 34.140000 0.490000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.130000 0.000000 29.270000 0.490000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.265000 0.000000 24.405000 0.490000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.400000 0.000000 19.540000 0.490000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.530000 0.000000 14.670000 0.490000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_ack_o
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.371 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.223 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 9.665000 0.000000 9.805000 0.490000 ;
    END
  END wbs_ack_o
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 481.765000 0.000000 481.905000 0.490000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 476.895000 0.000000 477.035000 0.490000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 472.030000 0.000000 472.170000 0.490000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 467.160000 0.000000 467.300000 0.490000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 462.295000 0.000000 462.435000 0.490000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 457.430000 0.000000 457.570000 0.490000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 452.560000 0.000000 452.700000 0.490000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 447.695000 0.000000 447.835000 0.490000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 442.825000 0.000000 442.965000 0.490000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 437.960000 0.000000 438.100000 0.490000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 433.095000 0.000000 433.235000 0.490000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 428.225000 0.000000 428.365000 0.490000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 423.360000 0.000000 423.500000 0.490000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 418.490000 0.000000 418.630000 0.490000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 413.625000 0.000000 413.765000 0.490000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 408.760000 0.000000 408.900000 0.490000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 403.890000 0.000000 404.030000 0.490000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 399.025000 0.000000 399.165000 0.490000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 394.155000 0.000000 394.295000 0.490000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 389.290000 0.000000 389.430000 0.490000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 384.425000 0.000000 384.565000 0.490000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 379.555000 0.000000 379.695000 0.490000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 374.690000 0.000000 374.830000 0.490000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 369.820000 0.000000 369.960000 0.490000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 364.955000 0.000000 365.095000 0.490000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 360.090000 0.000000 360.230000 0.490000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 355.220000 0.000000 355.360000 0.490000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 350.355000 0.000000 350.495000 0.490000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 345.485000 0.000000 345.625000 0.490000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 340.620000 0.000000 340.760000 0.490000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 335.755000 0.000000 335.895000 0.490000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 8.3682 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 41.209 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.7274 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 32.424 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met2 ;
        RECT 330.885000 0.000000 331.025000 0.490000 ;
    END
  END wbs_dat_o[0]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.940000 0.000000 1134.080000 0.490000 ;
    END
  END la_data_in[127]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1129.075000 0.000000 1129.215000 0.490000 ;
    END
  END la_data_in[126]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1124.205000 0.000000 1124.345000 0.490000 ;
    END
  END la_data_in[125]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.340000 0.000000 1119.480000 0.490000 ;
    END
  END la_data_in[124]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.475000 0.000000 1114.615000 0.490000 ;
    END
  END la_data_in[123]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.605000 0.000000 1109.745000 0.490000 ;
    END
  END la_data_in[122]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1104.740000 0.000000 1104.880000 0.490000 ;
    END
  END la_data_in[121]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1099.870000 0.000000 1100.010000 0.490000 ;
    END
  END la_data_in[120]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.005000 0.000000 1095.145000 0.490000 ;
    END
  END la_data_in[119]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.140000 0.000000 1090.280000 0.490000 ;
    END
  END la_data_in[118]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1085.270000 0.000000 1085.410000 0.490000 ;
    END
  END la_data_in[117]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.405000 0.000000 1080.545000 0.490000 ;
    END
  END la_data_in[116]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.535000 0.000000 1075.675000 0.490000 ;
    END
  END la_data_in[115]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.670000 0.000000 1070.810000 0.490000 ;
    END
  END la_data_in[114]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1065.805000 0.000000 1065.945000 0.490000 ;
    END
  END la_data_in[113]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.935000 0.000000 1061.075000 0.490000 ;
    END
  END la_data_in[112]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.070000 0.000000 1056.210000 0.490000 ;
    END
  END la_data_in[111]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1051.200000 0.000000 1051.340000 0.490000 ;
    END
  END la_data_in[110]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1046.335000 0.000000 1046.475000 0.490000 ;
    END
  END la_data_in[109]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1041.470000 0.000000 1041.610000 0.490000 ;
    END
  END la_data_in[108]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.600000 0.000000 1036.740000 0.490000 ;
    END
  END la_data_in[107]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.735000 0.000000 1031.875000 0.490000 ;
    END
  END la_data_in[106]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.865000 0.000000 1027.005000 0.490000 ;
    END
  END la_data_in[105]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.000000 0.000000 1022.140000 0.490000 ;
    END
  END la_data_in[104]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.135000 0.000000 1017.275000 0.490000 ;
    END
  END la_data_in[103]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1012.265000 0.000000 1012.405000 0.490000 ;
    END
  END la_data_in[102]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.400000 0.000000 1007.540000 0.490000 ;
    END
  END la_data_in[101]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1002.530000 0.000000 1002.670000 0.490000 ;
    END
  END la_data_in[100]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 997.665000 0.000000 997.805000 0.490000 ;
    END
  END la_data_in[99]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.800000 0.000000 992.940000 0.490000 ;
    END
  END la_data_in[98]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.930000 0.000000 988.070000 0.490000 ;
    END
  END la_data_in[97]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.065000 0.000000 983.205000 0.490000 ;
    END
  END la_data_in[96]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.195000 0.000000 978.335000 0.490000 ;
    END
  END la_data_in[95]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.330000 0.000000 973.470000 0.490000 ;
    END
  END la_data_in[94]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 968.465000 0.000000 968.605000 0.490000 ;
    END
  END la_data_in[93]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 963.595000 0.000000 963.735000 0.490000 ;
    END
  END la_data_in[92]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 958.730000 0.000000 958.870000 0.490000 ;
    END
  END la_data_in[91]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.860000 0.000000 954.000000 0.490000 ;
    END
  END la_data_in[90]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.995000 0.000000 949.135000 0.490000 ;
    END
  END la_data_in[89]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 944.130000 0.000000 944.270000 0.490000 ;
    END
  END la_data_in[88]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 939.260000 0.000000 939.400000 0.490000 ;
    END
  END la_data_in[87]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.395000 0.000000 934.535000 0.490000 ;
    END
  END la_data_in[86]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.525000 0.000000 929.665000 0.490000 ;
    END
  END la_data_in[85]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.660000 0.000000 924.800000 0.490000 ;
    END
  END la_data_in[84]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 919.795000 0.000000 919.935000 0.490000 ;
    END
  END la_data_in[83]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 914.925000 0.000000 915.065000 0.490000 ;
    END
  END la_data_in[82]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.060000 0.000000 910.200000 0.490000 ;
    END
  END la_data_in[81]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 905.190000 0.000000 905.330000 0.490000 ;
    END
  END la_data_in[80]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 900.325000 0.000000 900.465000 0.490000 ;
    END
  END la_data_in[79]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.460000 0.000000 895.600000 0.490000 ;
    END
  END la_data_in[78]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.590000 0.000000 890.730000 0.490000 ;
    END
  END la_data_in[77]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 885.725000 0.000000 885.865000 0.490000 ;
    END
  END la_data_in[76]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 880.855000 0.000000 880.995000 0.490000 ;
    END
  END la_data_in[75]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 875.990000 0.000000 876.130000 0.490000 ;
    END
  END la_data_in[74]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.125000 0.000000 871.265000 0.490000 ;
    END
  END la_data_in[73]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.255000 0.000000 866.395000 0.490000 ;
    END
  END la_data_in[72]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.390000 0.000000 861.530000 0.490000 ;
    END
  END la_data_in[71]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 856.520000 0.000000 856.660000 0.490000 ;
    END
  END la_data_in[70]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.655000 0.000000 851.795000 0.490000 ;
    END
  END la_data_in[69]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.790000 0.000000 846.930000 0.490000 ;
    END
  END la_data_in[68]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.920000 0.000000 842.060000 0.490000 ;
    END
  END la_data_in[67]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.055000 0.000000 837.195000 0.490000 ;
    END
  END la_data_in[66]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.185000 0.000000 832.325000 0.490000 ;
    END
  END la_data_in[65]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.320000 0.000000 827.460000 0.490000 ;
    END
  END la_data_in[64]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 822.455000 0.000000 822.595000 0.490000 ;
    END
  END la_data_in[63]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.585000 0.000000 817.725000 0.490000 ;
    END
  END la_data_in[62]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.720000 0.000000 812.860000 0.490000 ;
    END
  END la_data_in[61]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.850000 0.000000 807.990000 0.490000 ;
    END
  END la_data_in[60]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.985000 0.000000 803.125000 0.490000 ;
    END
  END la_data_in[59]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 798.120000 0.000000 798.260000 0.490000 ;
    END
  END la_data_in[58]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.250000 0.000000 793.390000 0.490000 ;
    END
  END la_data_in[57]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.385000 0.000000 788.525000 0.490000 ;
    END
  END la_data_in[56]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.515000 0.000000 783.655000 0.490000 ;
    END
  END la_data_in[55]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 778.650000 0.000000 778.790000 0.490000 ;
    END
  END la_data_in[54]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.785000 0.000000 773.925000 0.490000 ;
    END
  END la_data_in[53]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.915000 0.000000 769.055000 0.490000 ;
    END
  END la_data_in[52]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.050000 0.000000 764.190000 0.490000 ;
    END
  END la_data_in[51]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.180000 0.000000 759.320000 0.490000 ;
    END
  END la_data_in[50]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.315000 0.000000 754.455000 0.490000 ;
    END
  END la_data_in[49]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.450000 0.000000 749.590000 0.490000 ;
    END
  END la_data_in[48]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.580000 0.000000 744.720000 0.490000 ;
    END
  END la_data_in[47]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.715000 0.000000 739.855000 0.490000 ;
    END
  END la_data_in[46]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.845000 0.000000 734.985000 0.490000 ;
    END
  END la_data_in[45]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.980000 0.000000 730.120000 0.490000 ;
    END
  END la_data_in[44]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.115000 0.000000 725.255000 0.490000 ;
    END
  END la_data_in[43]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.245000 0.000000 720.385000 0.490000 ;
    END
  END la_data_in[42]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 715.380000 0.000000 715.520000 0.490000 ;
    END
  END la_data_in[41]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.510000 0.000000 710.650000 0.490000 ;
    END
  END la_data_in[40]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.645000 0.000000 705.785000 0.490000 ;
    END
  END la_data_in[39]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.780000 0.000000 700.920000 0.490000 ;
    END
  END la_data_in[38]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.910000 0.000000 696.050000 0.490000 ;
    END
  END la_data_in[37]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.045000 0.000000 691.185000 0.490000 ;
    END
  END la_data_in[36]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.175000 0.000000 686.315000 0.490000 ;
    END
  END la_data_in[35]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.310000 0.000000 681.450000 0.490000 ;
    END
  END la_data_in[34]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.445000 0.000000 676.585000 0.490000 ;
    END
  END la_data_in[33]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 671.575000 0.000000 671.715000 0.490000 ;
    END
  END la_data_in[32]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.710000 0.000000 666.850000 0.490000 ;
    END
  END la_data_in[31]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.840000 0.000000 661.980000 0.490000 ;
    END
  END la_data_in[30]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.975000 0.000000 657.115000 0.490000 ;
    END
  END la_data_in[29]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.110000 0.000000 652.250000 0.490000 ;
    END
  END la_data_in[28]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.240000 0.000000 647.380000 0.490000 ;
    END
  END la_data_in[27]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.375000 0.000000 642.515000 0.490000 ;
    END
  END la_data_in[26]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.505000 0.000000 637.645000 0.490000 ;
    END
  END la_data_in[25]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.640000 0.000000 632.780000 0.490000 ;
    END
  END la_data_in[24]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 627.775000 0.000000 627.915000 0.490000 ;
    END
  END la_data_in[23]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.905000 0.000000 623.045000 0.490000 ;
    END
  END la_data_in[22]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 618.040000 0.000000 618.180000 0.490000 ;
    END
  END la_data_in[21]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 613.170000 0.000000 613.310000 0.490000 ;
    END
  END la_data_in[20]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.305000 0.000000 608.445000 0.490000 ;
    END
  END la_data_in[19]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.440000 0.000000 603.580000 0.490000 ;
    END
  END la_data_in[18]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.570000 0.000000 598.710000 0.490000 ;
    END
  END la_data_in[17]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.705000 0.000000 593.845000 0.490000 ;
    END
  END la_data_in[16]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6552 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.158 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 588.835000 0.000000 588.975000 0.490000 ;
    END
  END la_data_in[15]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6566 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.165 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 583.970000 0.000000 584.110000 0.490000 ;
    END
  END la_data_in[14]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7693 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.728 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 579.105000 0.000000 579.245000 0.490000 ;
    END
  END la_data_in[13]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.8071 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.918 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 574.235000 0.000000 574.375000 0.490000 ;
    END
  END la_data_in[12]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6734 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.249 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 569.370000 0.000000 569.510000 0.490000 ;
    END
  END la_data_in[11]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.658 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.172 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 564.500000 0.000000 564.640000 0.490000 ;
    END
  END la_data_in[10]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6629 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.197 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 559.635000 0.000000 559.775000 0.490000 ;
    END
  END la_data_in[9]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7154 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.459 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 554.770000 0.000000 554.910000 0.490000 ;
    END
  END la_data_in[8]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.382 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 549.900000 0.000000 550.040000 0.490000 ;
    END
  END la_data_in[7]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6783 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.273 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 545.035000 0.000000 545.175000 0.490000 ;
    END
  END la_data_in[6]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7637 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.701 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 540.165000 0.000000 540.305000 0.490000 ;
    END
  END la_data_in[5]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7952 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.858 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 535.300000 0.000000 535.440000 0.490000 ;
    END
  END la_data_in[4]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7329 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.547 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 530.435000 0.000000 530.575000 0.490000 ;
    END
  END la_data_in[3]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7063 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.414 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 525.565000 0.000000 525.705000 0.490000 ;
    END
  END la_data_in[2]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.6958 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.361 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 520.700000 0.000000 520.840000 0.490000 ;
    END
  END la_data_in[1]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 52.7168 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 263.466 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 515.830000 0.000000 515.970000 0.490000 ;
    END
  END la_data_in[0]
  PIN la_data_out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1756.915000 0.000000 1757.055000 0.490000 ;
    END
  END la_data_out[127]
  PIN la_data_out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1752.050000 0.000000 1752.190000 0.490000 ;
    END
  END la_data_out[126]
  PIN la_data_out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1747.185000 0.000000 1747.325000 0.490000 ;
    END
  END la_data_out[125]
  PIN la_data_out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1742.315000 0.000000 1742.455000 0.490000 ;
    END
  END la_data_out[124]
  PIN la_data_out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1737.450000 0.000000 1737.590000 0.490000 ;
    END
  END la_data_out[123]
  PIN la_data_out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1732.580000 0.000000 1732.720000 0.490000 ;
    END
  END la_data_out[122]
  PIN la_data_out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1727.715000 0.000000 1727.855000 0.490000 ;
    END
  END la_data_out[121]
  PIN la_data_out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1722.850000 0.000000 1722.990000 0.490000 ;
    END
  END la_data_out[120]
  PIN la_data_out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1717.980000 0.000000 1718.120000 0.490000 ;
    END
  END la_data_out[119]
  PIN la_data_out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1713.115000 0.000000 1713.255000 0.490000 ;
    END
  END la_data_out[118]
  PIN la_data_out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1708.245000 0.000000 1708.385000 0.490000 ;
    END
  END la_data_out[117]
  PIN la_data_out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1703.380000 0.000000 1703.520000 0.490000 ;
    END
  END la_data_out[116]
  PIN la_data_out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1698.515000 0.000000 1698.655000 0.490000 ;
    END
  END la_data_out[115]
  PIN la_data_out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1693.645000 0.000000 1693.785000 0.490000 ;
    END
  END la_data_out[114]
  PIN la_data_out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1688.780000 0.000000 1688.920000 0.490000 ;
    END
  END la_data_out[113]
  PIN la_data_out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1683.910000 0.000000 1684.050000 0.490000 ;
    END
  END la_data_out[112]
  PIN la_data_out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1679.045000 0.000000 1679.185000 0.490000 ;
    END
  END la_data_out[111]
  PIN la_data_out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1674.180000 0.000000 1674.320000 0.490000 ;
    END
  END la_data_out[110]
  PIN la_data_out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1669.310000 0.000000 1669.450000 0.490000 ;
    END
  END la_data_out[109]
  PIN la_data_out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1664.445000 0.000000 1664.585000 0.490000 ;
    END
  END la_data_out[108]
  PIN la_data_out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1659.575000 0.000000 1659.715000 0.490000 ;
    END
  END la_data_out[107]
  PIN la_data_out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1654.710000 0.000000 1654.850000 0.490000 ;
    END
  END la_data_out[106]
  PIN la_data_out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1649.845000 0.000000 1649.985000 0.490000 ;
    END
  END la_data_out[105]
  PIN la_data_out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1644.975000 0.000000 1645.115000 0.490000 ;
    END
  END la_data_out[104]
  PIN la_data_out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1640.110000 0.000000 1640.250000 0.490000 ;
    END
  END la_data_out[103]
  PIN la_data_out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1635.240000 0.000000 1635.380000 0.490000 ;
    END
  END la_data_out[102]
  PIN la_data_out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1630.375000 0.000000 1630.515000 0.490000 ;
    END
  END la_data_out[101]
  PIN la_data_out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1625.510000 0.000000 1625.650000 0.490000 ;
    END
  END la_data_out[100]
  PIN la_data_out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1620.640000 0.000000 1620.780000 0.490000 ;
    END
  END la_data_out[99]
  PIN la_data_out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 140.755 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 652.804 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 594.303 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3105.49 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.46514 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1615.775000 0.000000 1615.915000 0.490000 ;
    END
  END la_data_out[98]
  PIN la_data_out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1610.905000 0.000000 1611.045000 0.490000 ;
    END
  END la_data_out[97]
  PIN la_data_out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1606.040000 0.000000 1606.180000 0.490000 ;
    END
  END la_data_out[96]
  PIN la_data_out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1601.175000 0.000000 1601.315000 0.490000 ;
    END
  END la_data_out[95]
  PIN la_data_out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1596.305000 0.000000 1596.445000 0.490000 ;
    END
  END la_data_out[94]
  PIN la_data_out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1591.440000 0.000000 1591.580000 0.490000 ;
    END
  END la_data_out[93]
  PIN la_data_out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1586.570000 0.000000 1586.710000 0.490000 ;
    END
  END la_data_out[92]
  PIN la_data_out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1581.705000 0.000000 1581.845000 0.490000 ;
    END
  END la_data_out[91]
  PIN la_data_out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.635 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.56 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.458 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 644.071 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 584.006 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.75 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1576.840000 0.000000 1576.980000 0.490000 ;
    END
  END la_data_out[90]
  PIN la_data_out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1571.970000 0.000000 1572.110000 0.490000 ;
    END
  END la_data_out[89]
  PIN la_data_out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1567.105000 0.000000 1567.245000 0.490000 ;
    END
  END la_data_out[88]
  PIN la_data_out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1562.235000 0.000000 1562.375000 0.490000 ;
    END
  END la_data_out[87]
  PIN la_data_out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1557.370000 0.000000 1557.510000 0.490000 ;
    END
  END la_data_out[86]
  PIN la_data_out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1552.505000 0.000000 1552.645000 0.490000 ;
    END
  END la_data_out[85]
  PIN la_data_out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1547.635000 0.000000 1547.775000 0.490000 ;
    END
  END la_data_out[84]
  PIN la_data_out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1542.770000 0.000000 1542.910000 0.490000 ;
    END
  END la_data_out[83]
  PIN la_data_out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1537.900000 0.000000 1538.040000 0.490000 ;
    END
  END la_data_out[82]
  PIN la_data_out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1533.035000 0.000000 1533.175000 0.490000 ;
    END
  END la_data_out[81]
  PIN la_data_out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1528.170000 0.000000 1528.310000 0.490000 ;
    END
  END la_data_out[80]
  PIN la_data_out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1523.300000 0.000000 1523.440000 0.490000 ;
    END
  END la_data_out[79]
  PIN la_data_out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1518.435000 0.000000 1518.575000 0.490000 ;
    END
  END la_data_out[78]
  PIN la_data_out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1513.565000 0.000000 1513.705000 0.490000 ;
    END
  END la_data_out[77]
  PIN la_data_out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1508.700000 0.000000 1508.840000 0.490000 ;
    END
  END la_data_out[76]
  PIN la_data_out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1503.835000 0.000000 1503.975000 0.490000 ;
    END
  END la_data_out[75]
  PIN la_data_out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 1498.965000 0.000000 1499.105000 0.490000 ;
    END
  END la_data_out[74]
  PIN la_data_out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.121 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 98.4503 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 483.366 LAYER met2  ;
    ANTENNAMAXCUTCAR 0.207677 LAYER via2  ;
    PORT
      LAYER met2 ;
        RECT 1494.100000 0.000000 1494.240000 0.490000 ;
    END
  END la_data_out[73]
  PIN la_data_out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1489.230000 0.000000 1489.370000 0.490000 ;
    END
  END la_data_out[72]
  PIN la_data_out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1484.365000 0.000000 1484.505000 0.490000 ;
    END
  END la_data_out[71]
  PIN la_data_out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1479.500000 0.000000 1479.640000 0.490000 ;
    END
  END la_data_out[70]
  PIN la_data_out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1474.630000 0.000000 1474.770000 0.490000 ;
    END
  END la_data_out[69]
  PIN la_data_out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1469.765000 0.000000 1469.905000 0.490000 ;
    END
  END la_data_out[68]
  PIN la_data_out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1464.895000 0.000000 1465.035000 0.490000 ;
    END
  END la_data_out[67]
  PIN la_data_out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1460.030000 0.000000 1460.170000 0.490000 ;
    END
  END la_data_out[66]
  PIN la_data_out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1455.165000 0.000000 1455.305000 0.490000 ;
    END
  END la_data_out[65]
  PIN la_data_out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1450.295000 0.000000 1450.435000 0.490000 ;
    END
  END la_data_out[64]
  PIN la_data_out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1445.430000 0.000000 1445.570000 0.490000 ;
    END
  END la_data_out[63]
  PIN la_data_out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1440.560000 0.000000 1440.700000 0.490000 ;
    END
  END la_data_out[62]
  PIN la_data_out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1435.695000 0.000000 1435.835000 0.490000 ;
    END
  END la_data_out[61]
  PIN la_data_out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1430.830000 0.000000 1430.970000 0.490000 ;
    END
  END la_data_out[60]
  PIN la_data_out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1425.960000 0.000000 1426.100000 0.490000 ;
    END
  END la_data_out[59]
  PIN la_data_out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1421.095000 0.000000 1421.235000 0.490000 ;
    END
  END la_data_out[58]
  PIN la_data_out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1416.225000 0.000000 1416.365000 0.490000 ;
    END
  END la_data_out[57]
  PIN la_data_out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1411.360000 0.000000 1411.500000 0.490000 ;
    END
  END la_data_out[56]
  PIN la_data_out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1406.495000 0.000000 1406.635000 0.490000 ;
    END
  END la_data_out[55]
  PIN la_data_out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1401.625000 0.000000 1401.765000 0.490000 ;
    END
  END la_data_out[54]
  PIN la_data_out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1396.760000 0.000000 1396.900000 0.490000 ;
    END
  END la_data_out[53]
  PIN la_data_out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1391.890000 0.000000 1392.030000 0.490000 ;
    END
  END la_data_out[52]
  PIN la_data_out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1387.025000 0.000000 1387.165000 0.490000 ;
    END
  END la_data_out[51]
  PIN la_data_out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1382.160000 0.000000 1382.300000 0.490000 ;
    END
  END la_data_out[50]
  PIN la_data_out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1377.290000 0.000000 1377.430000 0.490000 ;
    END
  END la_data_out[49]
  PIN la_data_out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1372.425000 0.000000 1372.565000 0.490000 ;
    END
  END la_data_out[48]
  PIN la_data_out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1367.555000 0.000000 1367.695000 0.490000 ;
    END
  END la_data_out[47]
  PIN la_data_out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1362.690000 0.000000 1362.830000 0.490000 ;
    END
  END la_data_out[46]
  PIN la_data_out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1357.825000 0.000000 1357.965000 0.490000 ;
    END
  END la_data_out[45]
  PIN la_data_out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1352.955000 0.000000 1353.095000 0.490000 ;
    END
  END la_data_out[44]
  PIN la_data_out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1348.090000 0.000000 1348.230000 0.490000 ;
    END
  END la_data_out[43]
  PIN la_data_out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1343.220000 0.000000 1343.360000 0.490000 ;
    END
  END la_data_out[42]
  PIN la_data_out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1338.355000 0.000000 1338.495000 0.490000 ;
    END
  END la_data_out[41]
  PIN la_data_out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1333.490000 0.000000 1333.630000 0.490000 ;
    END
  END la_data_out[40]
  PIN la_data_out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1328.620000 0.000000 1328.760000 0.490000 ;
    END
  END la_data_out[39]
  PIN la_data_out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1323.755000 0.000000 1323.895000 0.490000 ;
    END
  END la_data_out[38]
  PIN la_data_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1318.885000 0.000000 1319.025000 0.490000 ;
    END
  END la_data_out[37]
  PIN la_data_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1314.020000 0.000000 1314.160000 0.490000 ;
    END
  END la_data_out[36]
  PIN la_data_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1309.155000 0.000000 1309.295000 0.490000 ;
    END
  END la_data_out[35]
  PIN la_data_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1304.285000 0.000000 1304.425000 0.490000 ;
    END
  END la_data_out[34]
  PIN la_data_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1299.420000 0.000000 1299.560000 0.490000 ;
    END
  END la_data_out[33]
  PIN la_data_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1294.550000 0.000000 1294.690000 0.490000 ;
    END
  END la_data_out[32]
  PIN la_data_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1289.685000 0.000000 1289.825000 0.490000 ;
    END
  END la_data_out[31]
  PIN la_data_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1284.820000 0.000000 1284.960000 0.490000 ;
    END
  END la_data_out[30]
  PIN la_data_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1279.950000 0.000000 1280.090000 0.490000 ;
    END
  END la_data_out[29]
  PIN la_data_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1275.085000 0.000000 1275.225000 0.490000 ;
    END
  END la_data_out[28]
  PIN la_data_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1270.215000 0.000000 1270.355000 0.490000 ;
    END
  END la_data_out[27]
  PIN la_data_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1265.350000 0.000000 1265.490000 0.490000 ;
    END
  END la_data_out[26]
  PIN la_data_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1260.485000 0.000000 1260.625000 0.490000 ;
    END
  END la_data_out[25]
  PIN la_data_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1255.615000 0.000000 1255.755000 0.490000 ;
    END
  END la_data_out[24]
  PIN la_data_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1250.750000 0.000000 1250.890000 0.490000 ;
    END
  END la_data_out[23]
  PIN la_data_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1245.880000 0.000000 1246.020000 0.490000 ;
    END
  END la_data_out[22]
  PIN la_data_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1241.015000 0.000000 1241.155000 0.490000 ;
    END
  END la_data_out[21]
  PIN la_data_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1236.150000 0.000000 1236.290000 0.490000 ;
    END
  END la_data_out[20]
  PIN la_data_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1231.280000 0.000000 1231.420000 0.490000 ;
    END
  END la_data_out[19]
  PIN la_data_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1226.415000 0.000000 1226.555000 0.490000 ;
    END
  END la_data_out[18]
  PIN la_data_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1221.545000 0.000000 1221.685000 0.490000 ;
    END
  END la_data_out[17]
  PIN la_data_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1216.680000 0.000000 1216.820000 0.490000 ;
    END
  END la_data_out[16]
  PIN la_data_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1211.815000 0.000000 1211.955000 0.490000 ;
    END
  END la_data_out[15]
  PIN la_data_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1206.945000 0.000000 1207.085000 0.490000 ;
    END
  END la_data_out[14]
  PIN la_data_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1202.080000 0.000000 1202.220000 0.490000 ;
    END
  END la_data_out[13]
  PIN la_data_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1197.210000 0.000000 1197.350000 0.490000 ;
    END
  END la_data_out[12]
  PIN la_data_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1192.345000 0.000000 1192.485000 0.490000 ;
    END
  END la_data_out[11]
  PIN la_data_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1187.480000 0.000000 1187.620000 0.490000 ;
    END
  END la_data_out[10]
  PIN la_data_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1182.610000 0.000000 1182.750000 0.490000 ;
    END
  END la_data_out[9]
  PIN la_data_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1177.745000 0.000000 1177.885000 0.490000 ;
    END
  END la_data_out[8]
  PIN la_data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1172.875000 0.000000 1173.015000 0.490000 ;
    END
  END la_data_out[7]
  PIN la_data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.8117 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.142 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.2089 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.343 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1168.010000 0.000000 1168.150000 0.490000 ;
    END
  END la_data_out[6]
  PIN la_data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1163.145000 0.000000 1163.285000 0.490000 ;
    END
  END la_data_out[5]
  PIN la_data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1158.275000 0.000000 1158.415000 0.490000 ;
    END
  END la_data_out[4]
  PIN la_data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.121 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.259 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1153.410000 0.000000 1153.550000 0.490000 ;
    END
  END la_data_out[3]
  PIN la_data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.069 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.046 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1148.540000 0.000000 1148.680000 0.490000 ;
    END
  END la_data_out[2]
  PIN la_data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.797 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.121 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1495 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 477.259 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1143.675000 0.000000 1143.815000 0.490000 ;
    END
  END la_data_out[1]
  PIN la_data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.3406 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.7872 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 118.02 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.2475 LAYER met2  ;
    ANTENNAMAXAREACAR 96.1099 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 476.848 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1138.810000 0.000000 1138.950000 0.490000 ;
    END
  END la_data_out[0]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2379.895000 0.000000 2380.035000 0.490000 ;
    END
  END la_oenb[127]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.025000 0.000000 2375.165000 0.490000 ;
    END
  END la_oenb[126]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2370.160000 0.000000 2370.300000 0.490000 ;
    END
  END la_oenb[125]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2365.290000 0.000000 2365.430000 0.490000 ;
    END
  END la_oenb[124]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2360.425000 0.000000 2360.565000 0.490000 ;
    END
  END la_oenb[123]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.560000 0.000000 2355.700000 0.490000 ;
    END
  END la_oenb[122]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.690000 0.000000 2350.830000 0.490000 ;
    END
  END la_oenb[121]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.825000 0.000000 2345.965000 0.490000 ;
    END
  END la_oenb[120]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2340.955000 0.000000 2341.095000 0.490000 ;
    END
  END la_oenb[119]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.090000 0.000000 2336.230000 0.490000 ;
    END
  END la_oenb[118]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.225000 0.000000 2331.365000 0.490000 ;
    END
  END la_oenb[117]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2326.355000 0.000000 2326.495000 0.490000 ;
    END
  END la_oenb[116]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2321.490000 0.000000 2321.630000 0.490000 ;
    END
  END la_oenb[115]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2316.620000 0.000000 2316.760000 0.490000 ;
    END
  END la_oenb[114]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.755000 0.000000 2311.895000 0.490000 ;
    END
  END la_oenb[113]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.890000 0.000000 2307.030000 0.490000 ;
    END
  END la_oenb[112]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2302.020000 0.000000 2302.160000 0.490000 ;
    END
  END la_oenb[111]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2297.155000 0.000000 2297.295000 0.490000 ;
    END
  END la_oenb[110]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.285000 0.000000 2292.425000 0.490000 ;
    END
  END la_oenb[109]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.420000 0.000000 2287.560000 0.490000 ;
    END
  END la_oenb[108]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2282.555000 0.000000 2282.695000 0.490000 ;
    END
  END la_oenb[107]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2277.685000 0.000000 2277.825000 0.490000 ;
    END
  END la_oenb[106]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.820000 0.000000 2272.960000 0.490000 ;
    END
  END la_oenb[105]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2267.950000 0.000000 2268.090000 0.490000 ;
    END
  END la_oenb[104]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2263.085000 0.000000 2263.225000 0.490000 ;
    END
  END la_oenb[103]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2258.220000 0.000000 2258.360000 0.490000 ;
    END
  END la_oenb[102]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.350000 0.000000 2253.490000 0.490000 ;
    END
  END la_oenb[101]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.485000 0.000000 2248.625000 0.490000 ;
    END
  END la_oenb[100]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2243.615000 0.000000 2243.755000 0.490000 ;
    END
  END la_oenb[99]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2238.750000 0.000000 2238.890000 0.490000 ;
    END
  END la_oenb[98]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2233.885000 0.000000 2234.025000 0.490000 ;
    END
  END la_oenb[97]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.015000 0.000000 2229.155000 0.490000 ;
    END
  END la_oenb[96]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.150000 0.000000 2224.290000 0.490000 ;
    END
  END la_oenb[95]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2219.280000 0.000000 2219.420000 0.490000 ;
    END
  END la_oenb[94]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2214.415000 0.000000 2214.555000 0.490000 ;
    END
  END la_oenb[93]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.550000 0.000000 2209.690000 0.490000 ;
    END
  END la_oenb[92]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.680000 0.000000 2204.820000 0.490000 ;
    END
  END la_oenb[91]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2199.815000 0.000000 2199.955000 0.490000 ;
    END
  END la_oenb[90]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2194.945000 0.000000 2195.085000 0.490000 ;
    END
  END la_oenb[89]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.080000 0.000000 2190.220000 0.490000 ;
    END
  END la_oenb[88]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.215000 0.000000 2185.355000 0.490000 ;
    END
  END la_oenb[87]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2180.345000 0.000000 2180.485000 0.490000 ;
    END
  END la_oenb[86]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2175.480000 0.000000 2175.620000 0.490000 ;
    END
  END la_oenb[85]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2170.610000 0.000000 2170.750000 0.490000 ;
    END
  END la_oenb[84]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.745000 0.000000 2165.885000 0.490000 ;
    END
  END la_oenb[83]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.880000 0.000000 2161.020000 0.490000 ;
    END
  END la_oenb[82]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2156.010000 0.000000 2156.150000 0.490000 ;
    END
  END la_oenb[81]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.145000 0.000000 2151.285000 0.490000 ;
    END
  END la_oenb[80]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.275000 0.000000 2146.415000 0.490000 ;
    END
  END la_oenb[79]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.410000 0.000000 2141.550000 0.490000 ;
    END
  END la_oenb[78]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.545000 0.000000 2136.685000 0.490000 ;
    END
  END la_oenb[77]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2131.675000 0.000000 2131.815000 0.490000 ;
    END
  END la_oenb[76]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.810000 0.000000 2126.950000 0.490000 ;
    END
  END la_oenb[75]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.940000 0.000000 2122.080000 0.490000 ;
    END
  END la_oenb[74]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2117.075000 0.000000 2117.215000 0.490000 ;
    END
  END la_oenb[73]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.210000 0.000000 2112.350000 0.490000 ;
    END
  END la_oenb[72]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.340000 0.000000 2107.480000 0.490000 ;
    END
  END la_oenb[71]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.475000 0.000000 2102.615000 0.490000 ;
    END
  END la_oenb[70]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.605000 0.000000 2097.745000 0.490000 ;
    END
  END la_oenb[69]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2092.740000 0.000000 2092.880000 0.490000 ;
    END
  END la_oenb[68]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2087.875000 0.000000 2088.015000 0.490000 ;
    END
  END la_oenb[67]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.005000 0.000000 2083.145000 0.490000 ;
    END
  END la_oenb[66]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2078.140000 0.000000 2078.280000 0.490000 ;
    END
  END la_oenb[65]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2073.270000 0.000000 2073.410000 0.490000 ;
    END
  END la_oenb[64]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.405000 0.000000 2068.545000 0.490000 ;
    END
  END la_oenb[63]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.540000 0.000000 2063.680000 0.490000 ;
    END
  END la_oenb[62]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.670000 0.000000 2058.810000 0.490000 ;
    END
  END la_oenb[61]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.805000 0.000000 2053.945000 0.490000 ;
    END
  END la_oenb[60]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2048.935000 0.000000 2049.075000 0.490000 ;
    END
  END la_oenb[59]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.070000 0.000000 2044.210000 0.490000 ;
    END
  END la_oenb[58]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2039.205000 0.000000 2039.345000 0.490000 ;
    END
  END la_oenb[57]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2034.335000 0.000000 2034.475000 0.490000 ;
    END
  END la_oenb[56]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.470000 0.000000 2029.610000 0.490000 ;
    END
  END la_oenb[55]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.600000 0.000000 2024.740000 0.490000 ;
    END
  END la_oenb[54]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.735000 0.000000 2019.875000 0.490000 ;
    END
  END la_oenb[53]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.870000 0.000000 2015.010000 0.490000 ;
    END
  END la_oenb[52]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2010.000000 0.000000 2010.140000 0.490000 ;
    END
  END la_oenb[51]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.135000 0.000000 2005.275000 0.490000 ;
    END
  END la_oenb[50]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.265000 0.000000 2000.405000 0.490000 ;
    END
  END la_oenb[49]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1995.400000 0.000000 1995.540000 0.490000 ;
    END
  END la_oenb[48]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1990.535000 0.000000 1990.675000 0.490000 ;
    END
  END la_oenb[47]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.665000 0.000000 1985.805000 0.490000 ;
    END
  END la_oenb[46]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.800000 0.000000 1980.940000 0.490000 ;
    END
  END la_oenb[45]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.930000 0.000000 1976.070000 0.490000 ;
    END
  END la_oenb[44]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.065000 0.000000 1971.205000 0.490000 ;
    END
  END la_oenb[43]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.200000 0.000000 1966.340000 0.490000 ;
    END
  END la_oenb[42]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.330000 0.000000 1961.470000 0.490000 ;
    END
  END la_oenb[41]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.465000 0.000000 1956.605000 0.490000 ;
    END
  END la_oenb[40]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1951.595000 0.000000 1951.735000 0.490000 ;
    END
  END la_oenb[39]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1946.730000 0.000000 1946.870000 0.490000 ;
    END
  END la_oenb[38]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.865000 0.000000 1942.005000 0.490000 ;
    END
  END la_oenb[37]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.995000 0.000000 1937.135000 0.490000 ;
    END
  END la_oenb[36]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1932.130000 0.000000 1932.270000 0.490000 ;
    END
  END la_oenb[35]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1927.260000 0.000000 1927.400000 0.490000 ;
    END
  END la_oenb[34]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.395000 0.000000 1922.535000 0.490000 ;
    END
  END la_oenb[33]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.530000 0.000000 1917.670000 0.490000 ;
    END
  END la_oenb[32]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1912.660000 0.000000 1912.800000 0.490000 ;
    END
  END la_oenb[31]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1907.795000 0.000000 1907.935000 0.490000 ;
    END
  END la_oenb[30]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1902.925000 0.000000 1903.065000 0.490000 ;
    END
  END la_oenb[29]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.060000 0.000000 1898.200000 0.490000 ;
    END
  END la_oenb[28]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1893.195000 0.000000 1893.335000 0.490000 ;
    END
  END la_oenb[27]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.325000 0.000000 1888.465000 0.490000 ;
    END
  END la_oenb[26]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1883.460000 0.000000 1883.600000 0.490000 ;
    END
  END la_oenb[25]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.590000 0.000000 1878.730000 0.490000 ;
    END
  END la_oenb[24]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.725000 0.000000 1873.865000 0.490000 ;
    END
  END la_oenb[23]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1868.860000 0.000000 1869.000000 0.490000 ;
    END
  END la_oenb[22]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1863.990000 0.000000 1864.130000 0.490000 ;
    END
  END la_oenb[21]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.125000 0.000000 1859.265000 0.490000 ;
    END
  END la_oenb[20]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.255000 0.000000 1854.395000 0.490000 ;
    END
  END la_oenb[19]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1849.390000 0.000000 1849.530000 0.490000 ;
    END
  END la_oenb[18]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1844.525000 0.000000 1844.665000 0.490000 ;
    END
  END la_oenb[17]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.655000 0.000000 1839.795000 0.490000 ;
    END
  END la_oenb[16]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.790000 0.000000 1834.930000 0.490000 ;
    END
  END la_oenb[15]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1829.920000 0.000000 1830.060000 0.490000 ;
    END
  END la_oenb[14]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1825.055000 0.000000 1825.195000 0.490000 ;
    END
  END la_oenb[13]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.190000 0.000000 1820.330000 0.490000 ;
    END
  END la_oenb[12]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.320000 0.000000 1815.460000 0.490000 ;
    END
  END la_oenb[11]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.455000 0.000000 1810.595000 0.490000 ;
    END
  END la_oenb[10]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.585000 0.000000 1805.725000 0.490000 ;
    END
  END la_oenb[9]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1800.720000 0.000000 1800.860000 0.490000 ;
    END
  END la_oenb[8]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.855000 0.000000 1795.995000 0.490000 ;
    END
  END la_oenb[7]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.985000 0.000000 1791.125000 0.490000 ;
    END
  END la_oenb[6]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1786.120000 0.000000 1786.260000 0.490000 ;
    END
  END la_oenb[5]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.250000 0.000000 1781.390000 0.490000 ;
    END
  END la_oenb[4]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.385000 0.000000 1776.525000 0.490000 ;
    END
  END la_oenb[3]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.520000 0.000000 1771.660000 0.490000 ;
    END
  END la_oenb[2]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1766.650000 0.000000 1766.790000 0.490000 ;
    END
  END la_oenb[1]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1761.785000 0.000000 1761.925000 0.490000 ;
    END
  END la_oenb[0]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 97.960000 0.800000 98.260000 ;
    END
  END io_in[37]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.8984 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.12 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 245.130000 0.800000 245.430000 ;
    END
  END io_in[36]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.808 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 392.300000 0.800000 392.600000 ;
    END
  END io_in[35]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 3.896 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 588.520000 0.800000 588.820000 ;
    END
  END io_in[34]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.3449 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 23.168 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 784.745000 0.800000 785.045000 ;
    END
  END io_in[33]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 980.970000 0.800000 981.270000 ;
    END
  END io_in[32]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1177.195000 0.800000 1177.495000 ;
    END
  END io_in[31]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1373.420000 0.800000 1373.720000 ;
    END
  END io_in[30]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 21.2814 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 113.496 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1569.640000 0.800000 1569.940000 ;
    END
  END io_in[29]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 33.2079 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 177.104 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1765.865000 0.800000 1766.165000 ;
    END
  END io_in[28]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.2654 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.744 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1962.090000 0.800000 1962.390000 ;
    END
  END io_in[27]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.2859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 33.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2158.315000 0.800000 2158.615000 ;
    END
  END io_in[26]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 20.9634 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 111.8 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2354.540000 0.800000 2354.840000 ;
    END
  END io_in[25]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2664 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.416 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2550.760000 0.800000 2551.060000 ;
    END
  END io_in[24]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1662 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.605 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 137.060000 2599.490000 137.200000 2599.980000 ;
    END
  END io_in[23]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0353 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.951 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 411.325000 2599.490000 411.465000 2599.980000 ;
    END
  END io_in[22]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1452 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.5 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 685.590000 2599.490000 685.730000 2599.980000 ;
    END
  END io_in[21]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0437 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.992 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 959.855000 2599.490000 959.995000 2599.980000 ;
    END
  END io_in[20]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1032 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.29 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1234.120000 2599.490000 1234.260000 2599.980000 ;
    END
  END io_in[19]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0892 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.22 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1508.380000 2599.490000 1508.520000 2599.980000 ;
    END
  END io_in[18]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0745 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.146 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1782.645000 2599.490000 1782.785000 2599.980000 ;
    END
  END io_in[17]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.9418 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 224.483 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2056.910000 2599.490000 2057.050000 2599.980000 ;
    END
  END io_in[16]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.175000 2599.490000 2331.315000 2599.980000 ;
    END
  END io_in[15]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2499.800000 2399.820000 2500.100000 ;
    END
  END io_in[14]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 14.0049 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 74.688 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2299.805000 2399.820000 2300.105000 ;
    END
  END io_in[13]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.9264 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 68.936 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2099.810000 2399.820000 2100.110000 ;
    END
  END io_in[12]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 13.5024 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 72.008 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1899.810000 2399.820000 1900.110000 ;
    END
  END io_in[11]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.2859 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 65.52 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1699.815000 2399.820000 1700.115000 ;
    END
  END io_in[10]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1499.820000 2399.820000 1500.120000 ;
    END
  END io_in[9]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1299.825000 2399.820000 1300.125000 ;
    END
  END io_in[8]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 30.5334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 162.84 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1099.830000 2399.820000 1100.130000 ;
    END
  END io_in[7]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 899.830000 2399.820000 900.130000 ;
    END
  END io_in[6]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1419 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.752 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 749.835000 2399.820000 750.135000 ;
    END
  END io_in[5]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 599.840000 2399.820000 600.140000 ;
    END
  END io_in[4]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 449.840000 2399.820000 450.140000 ;
    END
  END io_in[3]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 12.4719 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 66.512 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 299.845000 2399.820000 300.145000 ;
    END
  END io_in[2]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 149.845000 2399.820000 150.145000 ;
    END
  END io_in[1]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 3.170000 2399.820000 3.470000 ;
    END
  END io_in[0]
  PIN io_out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5774 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.896 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 48.905000 0.800000 49.205000 ;
    END
  END io_out[37]
  PIN io_out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.6949 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.368 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 196.075000 0.800000 196.375000 ;
    END
  END io_out[36]
  PIN io_out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.8204 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 343.240000 0.800000 343.540000 ;
    END
  END io_out[35]
  PIN io_out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 11.9037 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 63.952 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 539.465000 0.800000 539.765000 ;
    END
  END io_out[34]
  PIN io_out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 10.9914 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 58.616 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 735.690000 0.800000 735.990000 ;
    END
  END io_out[33]
  PIN io_out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.2989 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 44.256 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 931.915000 0.800000 932.215000 ;
    END
  END io_out[32]
  PIN io_out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.7674 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 4.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1128.140000 0.800000 1128.440000 ;
    END
  END io_out[31]
  PIN io_out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.1334 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 38.04 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1324.360000 0.800000 1324.660000 ;
    END
  END io_out[30]
  PIN io_out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3009 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1520.585000 0.800000 1520.885000 ;
    END
  END io_out[29]
  PIN io_out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.4644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 34.472 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1716.810000 0.800000 1717.110000 ;
    END
  END io_out[28]
  PIN io_out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 7.5099 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 40.048 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1913.035000 0.800000 1913.335000 ;
    END
  END io_out[27]
  PIN io_out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 8.1864 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 43.656 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2109.260000 0.800000 2109.560000 ;
    END
  END io_out[26]
  PIN io_out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 6.8844 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 36.712 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2305.480000 0.800000 2305.780000 ;
    END
  END io_out[25]
  PIN io_out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.3729 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.984 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2501.705000 0.800000 2502.005000 ;
    END
  END io_out[24]
  PIN io_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1011 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.28 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 68.495000 2599.490000 68.635000 2599.980000 ;
    END
  END io_out[23]
  PIN io_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 43.9436 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.492 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 342.760000 2599.490000 342.900000 2599.980000 ;
    END
  END io_out[22]
  PIN io_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1417 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.482 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 617.025000 2599.490000 617.165000 2599.980000 ;
    END
  END io_out[21]
  PIN io_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0402 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.975 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 891.290000 2599.490000 891.430000 2599.980000 ;
    END
  END io_out[20]
  PIN io_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0542 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.045 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1165.550000 2599.490000 1165.690000 2599.980000 ;
    END
  END io_out[19]
  PIN io_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1613 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.58 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1439.815000 2599.490000 1439.955000 2599.980000 ;
    END
  END io_out[18]
  PIN io_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0304 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 219.926 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1714.080000 2599.490000 1714.220000 2599.980000 ;
    END
  END io_out[17]
  PIN io_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.0815 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.182 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1988.345000 2599.490000 1988.485000 2599.980000 ;
    END
  END io_out[16]
  PIN io_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 44.1648 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 220.598 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2262.610000 2599.490000 2262.750000 2599.980000 ;
    END
  END io_out[15]
  PIN io_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 18.1134 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 96.6 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2549.800000 2399.820000 2550.100000 ;
    END
  END io_out[14]
  PIN io_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2349.805000 2399.820000 2350.105000 ;
    END
  END io_out[13]
  PIN io_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.9272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 480.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2447.39 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2149.805000 2399.820000 2150.105000 ;
    END
  END io_out[12]
  PIN io_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.9272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 480.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2447.39 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1949.810000 2399.820000 1950.110000 ;
    END
  END io_out[11]
  PIN io_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1749.815000 2399.820000 1750.115000 ;
    END
  END io_out[10]
  PIN io_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2904 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.544 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1549.820000 2399.820000 1550.120000 ;
    END
  END io_out[9]
  PIN io_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.9799 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.888 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1349.825000 2399.820000 1350.125000 ;
    END
  END io_out[8]
  PIN io_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1149.825000 2399.820000 1150.125000 ;
    END
  END io_out[7]
  PIN io_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 4.5114 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 24.056 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 949.830000 2399.820000 950.130000 ;
    END
  END io_out[6]
  PIN io_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 799.835000 2399.820000 800.135000 ;
    END
  END io_out[5]
  PIN io_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.0589 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 26.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 649.835000 2399.820000 650.135000 ;
    END
  END io_out[4]
  PIN io_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 17.5584 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 93.64 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 499.840000 2399.820000 500.140000 ;
    END
  END io_out[3]
  PIN io_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.9272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 480.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2447.39 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 349.845000 2399.820000 350.145000 ;
    END
  END io_out[2]
  PIN io_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.1459 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 27.44 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 199.845000 2399.820000 200.145000 ;
    END
  END io_out[1]
  PIN io_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 5.6424 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 30.088 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 49.850000 2399.820000 50.150000 ;
    END
  END io_out[0]
  PIN io_oeb[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.608 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 1.460000 0.000000 1.760000 0.800000 ;
    END
  END io_oeb[37]
  PIN io_oeb[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 147.020000 0.800000 147.320000 ;
    END
  END io_oeb[36]
  PIN io_oeb[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.1644 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 0.872 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 294.185000 0.800000 294.485000 ;
    END
  END io_oeb[35]
  PIN io_oeb[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 7.9374 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 42.328 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 490.410000 0.800000 490.710000 ;
    END
  END io_oeb[34]
  PIN io_oeb[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 14.9169 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 79.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 686.635000 0.800000 686.935000 ;
    END
  END io_oeb[33]
  PIN io_oeb[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 882.860000 0.800000 883.160000 ;
    END
  END io_oeb[32]
  PIN io_oeb[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.891 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 5.5324 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 31.384 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1079.080000 0.800000 1079.380000 ;
    END
  END io_oeb[31]
  PIN io_oeb[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.2386 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 1.264 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNADIFFAREA 0.891 LAYER met4  ;
    ANTENNAPARTIALMETALAREA 59.1783 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 316.088 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1275.305000 0.800000 1275.605000 ;
    END
  END io_oeb[30]
  PIN io_oeb[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 32.6214 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 173.976 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1471.530000 0.800000 1471.830000 ;
    END
  END io_oeb[29]
  PIN io_oeb[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.6599 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.848 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1667.755000 0.800000 1668.055000 ;
    END
  END io_oeb[28]
  PIN io_oeb[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 28.8234 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 153.72 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1863.980000 0.800000 1864.280000 ;
    END
  END io_oeb[27]
  PIN io_oeb[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 24.2544 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 129.352 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2060.200000 0.800000 2060.500000 ;
    END
  END io_oeb[26]
  PIN io_oeb[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 20.3829 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 108.704 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2256.425000 0.800000 2256.725000 ;
    END
  END io_oeb[25]
  PIN io_oeb[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4455 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 0.4314 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 2.296 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2452.650000 0.800000 2452.950000 ;
    END
  END io_oeb[24]
  PIN io_oeb[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 19.5591 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 97.5695 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 2.460000 2599.495000 2.600000 2599.980000 ;
    END
  END io_oeb[23]
  PIN io_oeb[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.0681 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 104.997 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 274.195000 2599.490000 274.335000 2599.980000 ;
    END
  END io_oeb[22]
  PIN io_oeb[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 20.9708 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 104.51 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 548.460000 2599.490000 548.600000 2599.980000 ;
    END
  END io_oeb[21]
  PIN io_oeb[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.6706 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 113.127 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 822.720000 2599.490000 822.860000 2599.980000 ;
    END
  END io_oeb[20]
  PIN io_oeb[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 21.8213 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 108.763 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1096.985000 2599.490000 1097.125000 2599.980000 ;
    END
  END io_oeb[19]
  PIN io_oeb[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 23.0474 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 115.129 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1371.250000 2599.490000 1371.390000 2599.980000 ;
    END
  END io_oeb[18]
  PIN io_oeb[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.5089 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 112.318 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1645.515000 2599.490000 1645.655000 2599.980000 ;
    END
  END io_oeb[17]
  PIN io_oeb[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 22.5124 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 112.336 LAYER met2  ;
    PORT
      LAYER met2 ;
        RECT 1919.780000 2599.490000 1919.920000 2599.980000 ;
    END
  END io_oeb[16]
  PIN io_oeb[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 0.1645 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 0.6615 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 453.548 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2452.68 LAYER met3  ;
    PORT
      LAYER met2 ;
        RECT 2194.040000 2599.490000 2194.180000 2599.980000 ;
    END
  END io_oeb[15]
  PIN io_oeb[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2599.330000 2399.820000 2599.630000 ;
    END
  END io_oeb[14]
  PIN io_oeb[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5813 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 15.184 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2399.800000 2399.820000 2400.100000 ;
    END
  END io_oeb[13]
  PIN io_oeb[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 2.5363 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 14.464 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2199.805000 2399.820000 2200.105000 ;
    END
  END io_oeb[12]
  PIN io_oeb[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7716 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.44 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1999.810000 2399.820000 2000.110000 ;
    END
  END io_oeb[11]
  PIN io_oeb[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 1.7971 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 9.576 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1799.815000 2399.820000 1800.115000 ;
    END
  END io_oeb[10]
  PIN io_oeb[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.5744 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 168.392 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1599.820000 2399.820000 1600.120000 ;
    END
  END io_oeb[9]
  PIN io_oeb[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 31.2294 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 166.552 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1399.820000 2399.820000 1400.120000 ;
    END
  END io_oeb[8]
  PIN io_oeb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1199.825000 2399.820000 1200.125000 ;
    END
  END io_oeb[7]
  PIN io_oeb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 999.830000 2399.820000 1000.130000 ;
    END
  END io_oeb[6]
  PIN io_oeb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5542 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.848 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 849.835000 2399.820000 850.135000 ;
    END
  END io_oeb[5]
  PIN io_oeb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 699.835000 2399.820000 700.135000 ;
    END
  END io_oeb[4]
  PIN io_oeb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.0022 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.312 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.937 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2449.43 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 549.840000 2399.820000 550.140000 ;
    END
  END io_oeb[3]
  PIN io_oeb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAPARTIALMETALAREA 3.5092 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 20.128 LAYER met3  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via3  ;
    ANTENNAPARTIALMETALAREA 175.636 LAYER met4  ;
    ANTENNAPARTIALMETALSIDEAREA 937.184 LAYER met4  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 399.840000 2399.820000 400.140000 ;
    END
  END io_oeb[2]
  PIN io_oeb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 27.4629 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 146.464 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 249.845000 2399.820000 250.145000 ;
    END
  END io_oeb[1]
  PIN io_oeb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 88.9272 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 480.912 LAYER met3  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 452.556 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 2447.39 LAYER met3  ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 99.850000 2399.820000 100.150000 ;
    END
  END io_oeb[0]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 441.355000 0.800000 441.655000 ;
    END
  END analog_io[28]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 637.580000 0.800000 637.880000 ;
    END
  END analog_io[27]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 833.800000 0.800000 834.100000 ;
    END
  END analog_io[26]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1030.025000 0.800000 1030.325000 ;
    END
  END analog_io[25]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1226.250000 0.800000 1226.550000 ;
    END
  END analog_io[24]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1422.475000 0.800000 1422.775000 ;
    END
  END analog_io[23]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1618.700000 0.800000 1619.000000 ;
    END
  END analog_io[22]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 1814.920000 0.800000 1815.220000 ;
    END
  END analog_io[21]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2011.145000 0.800000 2011.445000 ;
    END
  END analog_io[20]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2207.370000 0.800000 2207.670000 ;
    END
  END analog_io[19]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2403.595000 0.800000 2403.895000 ;
    END
  END analog_io[18]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000000 2598.110000 0.800000 2598.410000 ;
    END
  END analog_io[17]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.630000 2599.490000 205.770000 2599.980000 ;
    END
  END analog_io[16]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.890000 2599.490000 480.030000 2599.980000 ;
    END
  END analog_io[15]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.155000 2599.490000 754.295000 2599.980000 ;
    END
  END analog_io[14]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.420000 2599.490000 1028.560000 2599.980000 ;
    END
  END analog_io[13]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.685000 2599.490000 1302.825000 2599.980000 ;
    END
  END analog_io[12]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1576.950000 2599.490000 1577.090000 2599.980000 ;
    END
  END analog_io[11]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1851.210000 2599.490000 1851.350000 2599.980000 ;
    END
  END analog_io[10]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2125.475000 2599.490000 2125.615000 2599.980000 ;
    END
  END analog_io[9]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2399.060000 2599.495000 2399.200000 2599.980000 ;
    END
  END analog_io[8]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2449.800000 2399.820000 2450.100000 ;
    END
  END analog_io[7]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2249.805000 2399.820000 2250.105000 ;
    END
  END analog_io[6]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 2049.810000 2399.820000 2050.110000 ;
    END
  END analog_io[5]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1849.815000 2399.820000 1850.115000 ;
    END
  END analog_io[4]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1649.815000 2399.820000 1650.115000 ;
    END
  END analog_io[3]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1449.820000 2399.820000 1450.120000 ;
    END
  END analog_io[2]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1249.825000 2399.820000 1250.125000 ;
    END
  END analog_io[1]
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2399.020000 1049.830000 2399.820000 1050.130000 ;
    END
  END analog_io[0]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.760000 0.000000 2384.900000 0.490000 ;
    END
  END user_clock2
  PIN user_irq[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2394.495000 0.000000 2394.635000 0.490000 ;
    END
  END user_irq[2]
  PIN user_irq[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6112 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.441 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.337 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.466 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.885 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.15 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2397.680000 0.000000 2397.820000 0.485000 ;
    END
  END user_irq[1]
  PIN user_irq[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4347 LAYER met2  ;
    ANTENNAPARTIALMETALAREA 25.6105 LAYER met2  ;
    ANTENNAPARTIALMETALSIDEAREA 126.437 LAYER met2  ;
    ANTENNAMODEL OXIDE1 ;
    ANTENNAGATEAREA 0.1965 LAYER met2  ;
    ANTENNAMAXAREACAR 130.333 LAYER met2  ;
    ANTENNAMAXSIDEAREACAR 643.448 LAYER met2  ;
    ANTENNAPARTIALCUTAREA 0.04 LAYER via2  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via2  ;
    ANTENNADIFFAREA 0.4347 LAYER met3  ;
    ANTENNAPARTIALMETALAREA 89.1222 LAYER met3  ;
    ANTENNAPARTIALMETALSIDEAREA 481.952 LAYER met3  ;
    ANTENNAGATEAREA 0.1965 LAYER met3  ;
    ANTENNAMAXAREACAR 583.881 LAYER met3  ;
    ANTENNAMAXSIDEAREACAR 3096.13 LAYER met3  ;
    ANTENNAMAXCUTCAR 0.203562 LAYER via3  ;
    PORT
      LAYER met2 ;
        RECT 2389.625000 0.000000 2389.765000 0.490000 ;
    END
  END user_irq[0]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2391.560000 6.260000 2393.300000 2592.000000 ;
    END
    PORT
      LAYER met4 ;
        RECT 6.520000 6.260000 8.320000 2592.020000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 750.655000 436.760000 752.395000 824.740000 ;
      LAYER met4 ;
        RECT 282.135000 436.760000 283.875000 824.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.655000 1367.760000 752.395000 1755.740000 ;
      LAYER met4 ;
        RECT 282.135000 1367.760000 283.875000 1755.740000 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.655000 1833.260000 752.395000 2221.240000 ;
      LAYER met4 ;
        RECT 282.135000 1833.260000 283.875000 2221.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.535000 431.220000 2179.275000 819.200000 ;
      LAYER met4 ;
        RECT 1709.015000 431.220000 1710.755000 819.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.535000 896.720000 2179.275000 1284.700000 ;
      LAYER met4 ;
        RECT 1709.015000 896.720000 1710.755000 1284.700000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.535000 1362.220000 2179.275000 1750.200000 ;
      LAYER met4 ;
        RECT 1709.015000 1362.220000 1710.755000 1750.200000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2177.535000 1827.720000 2179.275000 2215.700000 ;
      LAYER met4 ;
        RECT 1709.015000 1827.720000 1710.755000 2215.700000 ;
    END
    PORT
      LAYER met4 ;
        RECT 750.655000 902.260000 752.395000 1290.240000 ;
      LAYER met4 ;
        RECT 282.135000 902.260000 283.875000 1290.240000 ;
    END
    PORT
      LAYER met4 ;
        RECT 238.275000 381.715000 240.075000 2268.435000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2223.515000 381.715000 2225.315000 2268.435000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2395.100000 2.660000 2396.900000 2595.620000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2.920000 2.660000 4.720000 2595.620000 ;
    END

# P/G pin shape extracted from block 'azadi_soc_top'
    PORT
      LAYER met4 ;
        RECT 278.735000 433.360000 280.475000 828.140000 ;
      LAYER met4 ;
        RECT 754.055000 433.360000 755.795000 828.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.735000 1364.360000 280.475000 1759.140000 ;
      LAYER met4 ;
        RECT 754.055000 1364.360000 755.795000 1759.140000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.735000 1829.860000 280.475000 2224.640000 ;
      LAYER met4 ;
        RECT 754.055000 1829.860000 755.795000 2224.640000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1705.615000 427.820000 1707.355000 822.600000 ;
      LAYER met4 ;
        RECT 2180.935000 427.820000 2182.675000 822.600000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1705.615000 893.320000 1707.355000 1288.100000 ;
      LAYER met4 ;
        RECT 2180.935000 893.320000 2182.675000 1288.100000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1705.615000 1358.820000 1707.355000 1753.600000 ;
      LAYER met4 ;
        RECT 2180.935000 1358.820000 2182.675000 1753.600000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1705.615000 1824.320000 1707.355000 2219.100000 ;
      LAYER met4 ;
        RECT 2180.935000 1824.320000 2182.675000 2219.100000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.735000 898.860000 280.475000 1293.640000 ;
      LAYER met4 ;
        RECT 754.055000 898.860000 755.795000 1293.640000 ;
    END
    PORT
      LAYER met4 ;
        RECT 234.675000 378.115000 236.475000 2272.035000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.115000 378.115000 2228.915000 2272.035000 ;
    END
# end of P/G pin shape extracted from block 'azadi_soc_top'

  END vssd1
  OBS
    LAYER li1 ;
      RECT 0.000000 0.000000 2399.820000 2599.980000 ;
    LAYER met1 ;
      RECT 0.000000 0.000000 2399.820000 2599.980000 ;
    LAYER met2 ;
      RECT 2399.340000 2599.355000 2399.820000 2599.980000 ;
      RECT 2331.455000 2599.355000 2398.920000 2599.980000 ;
      RECT 2.740000 2599.355000 68.355000 2599.980000 ;
      RECT 0.000000 2599.355000 2.320000 2599.980000 ;
      RECT 2331.455000 2599.350000 2399.820000 2599.355000 ;
      RECT 2262.890000 2599.350000 2331.035000 2599.980000 ;
      RECT 2194.320000 2599.350000 2262.470000 2599.980000 ;
      RECT 2125.755000 2599.350000 2193.900000 2599.980000 ;
      RECT 2057.190000 2599.350000 2125.335000 2599.980000 ;
      RECT 1988.625000 2599.350000 2056.770000 2599.980000 ;
      RECT 1920.060000 2599.350000 1988.205000 2599.980000 ;
      RECT 1851.490000 2599.350000 1919.640000 2599.980000 ;
      RECT 1782.925000 2599.350000 1851.070000 2599.980000 ;
      RECT 1714.360000 2599.350000 1782.505000 2599.980000 ;
      RECT 1645.795000 2599.350000 1713.940000 2599.980000 ;
      RECT 1577.230000 2599.350000 1645.375000 2599.980000 ;
      RECT 1508.660000 2599.350000 1576.810000 2599.980000 ;
      RECT 1440.095000 2599.350000 1508.240000 2599.980000 ;
      RECT 1371.530000 2599.350000 1439.675000 2599.980000 ;
      RECT 1302.965000 2599.350000 1371.110000 2599.980000 ;
      RECT 1234.400000 2599.350000 1302.545000 2599.980000 ;
      RECT 1165.830000 2599.350000 1233.980000 2599.980000 ;
      RECT 1097.265000 2599.350000 1165.410000 2599.980000 ;
      RECT 1028.700000 2599.350000 1096.845000 2599.980000 ;
      RECT 960.135000 2599.350000 1028.280000 2599.980000 ;
      RECT 891.570000 2599.350000 959.715000 2599.980000 ;
      RECT 823.000000 2599.350000 891.150000 2599.980000 ;
      RECT 754.435000 2599.350000 822.580000 2599.980000 ;
      RECT 685.870000 2599.350000 754.015000 2599.980000 ;
      RECT 617.305000 2599.350000 685.450000 2599.980000 ;
      RECT 548.740000 2599.350000 616.885000 2599.980000 ;
      RECT 480.170000 2599.350000 548.320000 2599.980000 ;
      RECT 411.605000 2599.350000 479.750000 2599.980000 ;
      RECT 343.040000 2599.350000 411.185000 2599.980000 ;
      RECT 274.475000 2599.350000 342.620000 2599.980000 ;
      RECT 205.910000 2599.350000 274.055000 2599.980000 ;
      RECT 137.340000 2599.350000 205.490000 2599.980000 ;
      RECT 68.775000 2599.350000 136.920000 2599.980000 ;
      RECT 0.000000 2599.350000 68.355000 2599.355000 ;
      RECT 0.000000 1.400000 2399.820000 2599.350000 ;
      RECT 0.625000 0.980000 2399.820000 1.400000 ;
      RECT 0.000000 0.630000 2399.820000 0.980000 ;
      RECT 2394.775000 0.625000 2399.820000 0.630000 ;
      RECT 2397.960000 0.000000 2399.820000 0.625000 ;
      RECT 2394.775000 0.000000 2397.540000 0.625000 ;
      RECT 2389.905000 0.000000 2394.355000 0.630000 ;
      RECT 2385.040000 0.000000 2389.485000 0.630000 ;
      RECT 2380.175000 0.000000 2384.620000 0.630000 ;
      RECT 2375.305000 0.000000 2379.755000 0.630000 ;
      RECT 2370.440000 0.000000 2374.885000 0.630000 ;
      RECT 2365.570000 0.000000 2370.020000 0.630000 ;
      RECT 2360.705000 0.000000 2365.150000 0.630000 ;
      RECT 2355.840000 0.000000 2360.285000 0.630000 ;
      RECT 2350.970000 0.000000 2355.420000 0.630000 ;
      RECT 2346.105000 0.000000 2350.550000 0.630000 ;
      RECT 2341.235000 0.000000 2345.685000 0.630000 ;
      RECT 2336.370000 0.000000 2340.815000 0.630000 ;
      RECT 2331.505000 0.000000 2335.950000 0.630000 ;
      RECT 2326.635000 0.000000 2331.085000 0.630000 ;
      RECT 2321.770000 0.000000 2326.215000 0.630000 ;
      RECT 2316.900000 0.000000 2321.350000 0.630000 ;
      RECT 2312.035000 0.000000 2316.480000 0.630000 ;
      RECT 2307.170000 0.000000 2311.615000 0.630000 ;
      RECT 2302.300000 0.000000 2306.750000 0.630000 ;
      RECT 2297.435000 0.000000 2301.880000 0.630000 ;
      RECT 2292.565000 0.000000 2297.015000 0.630000 ;
      RECT 2287.700000 0.000000 2292.145000 0.630000 ;
      RECT 2282.835000 0.000000 2287.280000 0.630000 ;
      RECT 2277.965000 0.000000 2282.415000 0.630000 ;
      RECT 2273.100000 0.000000 2277.545000 0.630000 ;
      RECT 2268.230000 0.000000 2272.680000 0.630000 ;
      RECT 2263.365000 0.000000 2267.810000 0.630000 ;
      RECT 2258.500000 0.000000 2262.945000 0.630000 ;
      RECT 2253.630000 0.000000 2258.080000 0.630000 ;
      RECT 2248.765000 0.000000 2253.210000 0.630000 ;
      RECT 2243.895000 0.000000 2248.345000 0.630000 ;
      RECT 2239.030000 0.000000 2243.475000 0.630000 ;
      RECT 2234.165000 0.000000 2238.610000 0.630000 ;
      RECT 2229.295000 0.000000 2233.745000 0.630000 ;
      RECT 2224.430000 0.000000 2228.875000 0.630000 ;
      RECT 2219.560000 0.000000 2224.010000 0.630000 ;
      RECT 2214.695000 0.000000 2219.140000 0.630000 ;
      RECT 2209.830000 0.000000 2214.275000 0.630000 ;
      RECT 2204.960000 0.000000 2209.410000 0.630000 ;
      RECT 2200.095000 0.000000 2204.540000 0.630000 ;
      RECT 2195.225000 0.000000 2199.675000 0.630000 ;
      RECT 2190.360000 0.000000 2194.805000 0.630000 ;
      RECT 2185.495000 0.000000 2189.940000 0.630000 ;
      RECT 2180.625000 0.000000 2185.075000 0.630000 ;
      RECT 2175.760000 0.000000 2180.205000 0.630000 ;
      RECT 2170.890000 0.000000 2175.340000 0.630000 ;
      RECT 2166.025000 0.000000 2170.470000 0.630000 ;
      RECT 2161.160000 0.000000 2165.605000 0.630000 ;
      RECT 2156.290000 0.000000 2160.740000 0.630000 ;
      RECT 2151.425000 0.000000 2155.870000 0.630000 ;
      RECT 2146.555000 0.000000 2151.005000 0.630000 ;
      RECT 2141.690000 0.000000 2146.135000 0.630000 ;
      RECT 2136.825000 0.000000 2141.270000 0.630000 ;
      RECT 2131.955000 0.000000 2136.405000 0.630000 ;
      RECT 2127.090000 0.000000 2131.535000 0.630000 ;
      RECT 2122.220000 0.000000 2126.670000 0.630000 ;
      RECT 2117.355000 0.000000 2121.800000 0.630000 ;
      RECT 2112.490000 0.000000 2116.935000 0.630000 ;
      RECT 2107.620000 0.000000 2112.070000 0.630000 ;
      RECT 2102.755000 0.000000 2107.200000 0.630000 ;
      RECT 2097.885000 0.000000 2102.335000 0.630000 ;
      RECT 2093.020000 0.000000 2097.465000 0.630000 ;
      RECT 2088.155000 0.000000 2092.600000 0.630000 ;
      RECT 2083.285000 0.000000 2087.735000 0.630000 ;
      RECT 2078.420000 0.000000 2082.865000 0.630000 ;
      RECT 2073.550000 0.000000 2078.000000 0.630000 ;
      RECT 2068.685000 0.000000 2073.130000 0.630000 ;
      RECT 2063.820000 0.000000 2068.265000 0.630000 ;
      RECT 2058.950000 0.000000 2063.400000 0.630000 ;
      RECT 2054.085000 0.000000 2058.530000 0.630000 ;
      RECT 2049.215000 0.000000 2053.665000 0.630000 ;
      RECT 2044.350000 0.000000 2048.795000 0.630000 ;
      RECT 2039.485000 0.000000 2043.930000 0.630000 ;
      RECT 2034.615000 0.000000 2039.065000 0.630000 ;
      RECT 2029.750000 0.000000 2034.195000 0.630000 ;
      RECT 2024.880000 0.000000 2029.330000 0.630000 ;
      RECT 2020.015000 0.000000 2024.460000 0.630000 ;
      RECT 2015.150000 0.000000 2019.595000 0.630000 ;
      RECT 2010.280000 0.000000 2014.730000 0.630000 ;
      RECT 2005.415000 0.000000 2009.860000 0.630000 ;
      RECT 2000.545000 0.000000 2004.995000 0.630000 ;
      RECT 1995.680000 0.000000 2000.125000 0.630000 ;
      RECT 1990.815000 0.000000 1995.260000 0.630000 ;
      RECT 1985.945000 0.000000 1990.395000 0.630000 ;
      RECT 1981.080000 0.000000 1985.525000 0.630000 ;
      RECT 1976.210000 0.000000 1980.660000 0.630000 ;
      RECT 1971.345000 0.000000 1975.790000 0.630000 ;
      RECT 1966.480000 0.000000 1970.925000 0.630000 ;
      RECT 1961.610000 0.000000 1966.060000 0.630000 ;
      RECT 1956.745000 0.000000 1961.190000 0.630000 ;
      RECT 1951.875000 0.000000 1956.325000 0.630000 ;
      RECT 1947.010000 0.000000 1951.455000 0.630000 ;
      RECT 1942.145000 0.000000 1946.590000 0.630000 ;
      RECT 1937.275000 0.000000 1941.725000 0.630000 ;
      RECT 1932.410000 0.000000 1936.855000 0.630000 ;
      RECT 1927.540000 0.000000 1931.990000 0.630000 ;
      RECT 1922.675000 0.000000 1927.120000 0.630000 ;
      RECT 1917.810000 0.000000 1922.255000 0.630000 ;
      RECT 1912.940000 0.000000 1917.390000 0.630000 ;
      RECT 1908.075000 0.000000 1912.520000 0.630000 ;
      RECT 1903.205000 0.000000 1907.655000 0.630000 ;
      RECT 1898.340000 0.000000 1902.785000 0.630000 ;
      RECT 1893.475000 0.000000 1897.920000 0.630000 ;
      RECT 1888.605000 0.000000 1893.055000 0.630000 ;
      RECT 1883.740000 0.000000 1888.185000 0.630000 ;
      RECT 1878.870000 0.000000 1883.320000 0.630000 ;
      RECT 1874.005000 0.000000 1878.450000 0.630000 ;
      RECT 1869.140000 0.000000 1873.585000 0.630000 ;
      RECT 1864.270000 0.000000 1868.720000 0.630000 ;
      RECT 1859.405000 0.000000 1863.850000 0.630000 ;
      RECT 1854.535000 0.000000 1858.985000 0.630000 ;
      RECT 1849.670000 0.000000 1854.115000 0.630000 ;
      RECT 1844.805000 0.000000 1849.250000 0.630000 ;
      RECT 1839.935000 0.000000 1844.385000 0.630000 ;
      RECT 1835.070000 0.000000 1839.515000 0.630000 ;
      RECT 1830.200000 0.000000 1834.650000 0.630000 ;
      RECT 1825.335000 0.000000 1829.780000 0.630000 ;
      RECT 1820.470000 0.000000 1824.915000 0.630000 ;
      RECT 1815.600000 0.000000 1820.050000 0.630000 ;
      RECT 1810.735000 0.000000 1815.180000 0.630000 ;
      RECT 1805.865000 0.000000 1810.315000 0.630000 ;
      RECT 1801.000000 0.000000 1805.445000 0.630000 ;
      RECT 1796.135000 0.000000 1800.580000 0.630000 ;
      RECT 1791.265000 0.000000 1795.715000 0.630000 ;
      RECT 1786.400000 0.000000 1790.845000 0.630000 ;
      RECT 1781.530000 0.000000 1785.980000 0.630000 ;
      RECT 1776.665000 0.000000 1781.110000 0.630000 ;
      RECT 1771.800000 0.000000 1776.245000 0.630000 ;
      RECT 1766.930000 0.000000 1771.380000 0.630000 ;
      RECT 1762.065000 0.000000 1766.510000 0.630000 ;
      RECT 1757.195000 0.000000 1761.645000 0.630000 ;
      RECT 1752.330000 0.000000 1756.775000 0.630000 ;
      RECT 1747.465000 0.000000 1751.910000 0.630000 ;
      RECT 1742.595000 0.000000 1747.045000 0.630000 ;
      RECT 1737.730000 0.000000 1742.175000 0.630000 ;
      RECT 1732.860000 0.000000 1737.310000 0.630000 ;
      RECT 1727.995000 0.000000 1732.440000 0.630000 ;
      RECT 1723.130000 0.000000 1727.575000 0.630000 ;
      RECT 1718.260000 0.000000 1722.710000 0.630000 ;
      RECT 1713.395000 0.000000 1717.840000 0.630000 ;
      RECT 1708.525000 0.000000 1712.975000 0.630000 ;
      RECT 1703.660000 0.000000 1708.105000 0.630000 ;
      RECT 1698.795000 0.000000 1703.240000 0.630000 ;
      RECT 1693.925000 0.000000 1698.375000 0.630000 ;
      RECT 1689.060000 0.000000 1693.505000 0.630000 ;
      RECT 1684.190000 0.000000 1688.640000 0.630000 ;
      RECT 1679.325000 0.000000 1683.770000 0.630000 ;
      RECT 1674.460000 0.000000 1678.905000 0.630000 ;
      RECT 1669.590000 0.000000 1674.040000 0.630000 ;
      RECT 1664.725000 0.000000 1669.170000 0.630000 ;
      RECT 1659.855000 0.000000 1664.305000 0.630000 ;
      RECT 1654.990000 0.000000 1659.435000 0.630000 ;
      RECT 1650.125000 0.000000 1654.570000 0.630000 ;
      RECT 1645.255000 0.000000 1649.705000 0.630000 ;
      RECT 1640.390000 0.000000 1644.835000 0.630000 ;
      RECT 1635.520000 0.000000 1639.970000 0.630000 ;
      RECT 1630.655000 0.000000 1635.100000 0.630000 ;
      RECT 1625.790000 0.000000 1630.235000 0.630000 ;
      RECT 1620.920000 0.000000 1625.370000 0.630000 ;
      RECT 1616.055000 0.000000 1620.500000 0.630000 ;
      RECT 1611.185000 0.000000 1615.635000 0.630000 ;
      RECT 1606.320000 0.000000 1610.765000 0.630000 ;
      RECT 1601.455000 0.000000 1605.900000 0.630000 ;
      RECT 1596.585000 0.000000 1601.035000 0.630000 ;
      RECT 1591.720000 0.000000 1596.165000 0.630000 ;
      RECT 1586.850000 0.000000 1591.300000 0.630000 ;
      RECT 1581.985000 0.000000 1586.430000 0.630000 ;
      RECT 1577.120000 0.000000 1581.565000 0.630000 ;
      RECT 1572.250000 0.000000 1576.700000 0.630000 ;
      RECT 1567.385000 0.000000 1571.830000 0.630000 ;
      RECT 1562.515000 0.000000 1566.965000 0.630000 ;
      RECT 1557.650000 0.000000 1562.095000 0.630000 ;
      RECT 1552.785000 0.000000 1557.230000 0.630000 ;
      RECT 1547.915000 0.000000 1552.365000 0.630000 ;
      RECT 1543.050000 0.000000 1547.495000 0.630000 ;
      RECT 1538.180000 0.000000 1542.630000 0.630000 ;
      RECT 1533.315000 0.000000 1537.760000 0.630000 ;
      RECT 1528.450000 0.000000 1532.895000 0.630000 ;
      RECT 1523.580000 0.000000 1528.030000 0.630000 ;
      RECT 1518.715000 0.000000 1523.160000 0.630000 ;
      RECT 1513.845000 0.000000 1518.295000 0.630000 ;
      RECT 1508.980000 0.000000 1513.425000 0.630000 ;
      RECT 1504.115000 0.000000 1508.560000 0.630000 ;
      RECT 1499.245000 0.000000 1503.695000 0.630000 ;
      RECT 1494.380000 0.000000 1498.825000 0.630000 ;
      RECT 1489.510000 0.000000 1493.960000 0.630000 ;
      RECT 1484.645000 0.000000 1489.090000 0.630000 ;
      RECT 1479.780000 0.000000 1484.225000 0.630000 ;
      RECT 1474.910000 0.000000 1479.360000 0.630000 ;
      RECT 1470.045000 0.000000 1474.490000 0.630000 ;
      RECT 1465.175000 0.000000 1469.625000 0.630000 ;
      RECT 1460.310000 0.000000 1464.755000 0.630000 ;
      RECT 1455.445000 0.000000 1459.890000 0.630000 ;
      RECT 1450.575000 0.000000 1455.025000 0.630000 ;
      RECT 1445.710000 0.000000 1450.155000 0.630000 ;
      RECT 1440.840000 0.000000 1445.290000 0.630000 ;
      RECT 1435.975000 0.000000 1440.420000 0.630000 ;
      RECT 1431.110000 0.000000 1435.555000 0.630000 ;
      RECT 1426.240000 0.000000 1430.690000 0.630000 ;
      RECT 1421.375000 0.000000 1425.820000 0.630000 ;
      RECT 1416.505000 0.000000 1420.955000 0.630000 ;
      RECT 1411.640000 0.000000 1416.085000 0.630000 ;
      RECT 1406.775000 0.000000 1411.220000 0.630000 ;
      RECT 1401.905000 0.000000 1406.355000 0.630000 ;
      RECT 1397.040000 0.000000 1401.485000 0.630000 ;
      RECT 1392.170000 0.000000 1396.620000 0.630000 ;
      RECT 1387.305000 0.000000 1391.750000 0.630000 ;
      RECT 1382.440000 0.000000 1386.885000 0.630000 ;
      RECT 1377.570000 0.000000 1382.020000 0.630000 ;
      RECT 1372.705000 0.000000 1377.150000 0.630000 ;
      RECT 1367.835000 0.000000 1372.285000 0.630000 ;
      RECT 1362.970000 0.000000 1367.415000 0.630000 ;
      RECT 1358.105000 0.000000 1362.550000 0.630000 ;
      RECT 1353.235000 0.000000 1357.685000 0.630000 ;
      RECT 1348.370000 0.000000 1352.815000 0.630000 ;
      RECT 1343.500000 0.000000 1347.950000 0.630000 ;
      RECT 1338.635000 0.000000 1343.080000 0.630000 ;
      RECT 1333.770000 0.000000 1338.215000 0.630000 ;
      RECT 1328.900000 0.000000 1333.350000 0.630000 ;
      RECT 1324.035000 0.000000 1328.480000 0.630000 ;
      RECT 1319.165000 0.000000 1323.615000 0.630000 ;
      RECT 1314.300000 0.000000 1318.745000 0.630000 ;
      RECT 1309.435000 0.000000 1313.880000 0.630000 ;
      RECT 1304.565000 0.000000 1309.015000 0.630000 ;
      RECT 1299.700000 0.000000 1304.145000 0.630000 ;
      RECT 1294.830000 0.000000 1299.280000 0.630000 ;
      RECT 1289.965000 0.000000 1294.410000 0.630000 ;
      RECT 1285.100000 0.000000 1289.545000 0.630000 ;
      RECT 1280.230000 0.000000 1284.680000 0.630000 ;
      RECT 1275.365000 0.000000 1279.810000 0.630000 ;
      RECT 1270.495000 0.000000 1274.945000 0.630000 ;
      RECT 1265.630000 0.000000 1270.075000 0.630000 ;
      RECT 1260.765000 0.000000 1265.210000 0.630000 ;
      RECT 1255.895000 0.000000 1260.345000 0.630000 ;
      RECT 1251.030000 0.000000 1255.475000 0.630000 ;
      RECT 1246.160000 0.000000 1250.610000 0.630000 ;
      RECT 1241.295000 0.000000 1245.740000 0.630000 ;
      RECT 1236.430000 0.000000 1240.875000 0.630000 ;
      RECT 1231.560000 0.000000 1236.010000 0.630000 ;
      RECT 1226.695000 0.000000 1231.140000 0.630000 ;
      RECT 1221.825000 0.000000 1226.275000 0.630000 ;
      RECT 1216.960000 0.000000 1221.405000 0.630000 ;
      RECT 1212.095000 0.000000 1216.540000 0.630000 ;
      RECT 1207.225000 0.000000 1211.675000 0.630000 ;
      RECT 1202.360000 0.000000 1206.805000 0.630000 ;
      RECT 1197.490000 0.000000 1201.940000 0.630000 ;
      RECT 1192.625000 0.000000 1197.070000 0.630000 ;
      RECT 1187.760000 0.000000 1192.205000 0.630000 ;
      RECT 1182.890000 0.000000 1187.340000 0.630000 ;
      RECT 1178.025000 0.000000 1182.470000 0.630000 ;
      RECT 1173.155000 0.000000 1177.605000 0.630000 ;
      RECT 1168.290000 0.000000 1172.735000 0.630000 ;
      RECT 1163.425000 0.000000 1167.870000 0.630000 ;
      RECT 1158.555000 0.000000 1163.005000 0.630000 ;
      RECT 1153.690000 0.000000 1158.135000 0.630000 ;
      RECT 1148.820000 0.000000 1153.270000 0.630000 ;
      RECT 1143.955000 0.000000 1148.400000 0.630000 ;
      RECT 1139.090000 0.000000 1143.535000 0.630000 ;
      RECT 1134.220000 0.000000 1138.670000 0.630000 ;
      RECT 1129.355000 0.000000 1133.800000 0.630000 ;
      RECT 1124.485000 0.000000 1128.935000 0.630000 ;
      RECT 1119.620000 0.000000 1124.065000 0.630000 ;
      RECT 1114.755000 0.000000 1119.200000 0.630000 ;
      RECT 1109.885000 0.000000 1114.335000 0.630000 ;
      RECT 1105.020000 0.000000 1109.465000 0.630000 ;
      RECT 1100.150000 0.000000 1104.600000 0.630000 ;
      RECT 1095.285000 0.000000 1099.730000 0.630000 ;
      RECT 1090.420000 0.000000 1094.865000 0.630000 ;
      RECT 1085.550000 0.000000 1090.000000 0.630000 ;
      RECT 1080.685000 0.000000 1085.130000 0.630000 ;
      RECT 1075.815000 0.000000 1080.265000 0.630000 ;
      RECT 1070.950000 0.000000 1075.395000 0.630000 ;
      RECT 1066.085000 0.000000 1070.530000 0.630000 ;
      RECT 1061.215000 0.000000 1065.665000 0.630000 ;
      RECT 1056.350000 0.000000 1060.795000 0.630000 ;
      RECT 1051.480000 0.000000 1055.930000 0.630000 ;
      RECT 1046.615000 0.000000 1051.060000 0.630000 ;
      RECT 1041.750000 0.000000 1046.195000 0.630000 ;
      RECT 1036.880000 0.000000 1041.330000 0.630000 ;
      RECT 1032.015000 0.000000 1036.460000 0.630000 ;
      RECT 1027.145000 0.000000 1031.595000 0.630000 ;
      RECT 1022.280000 0.000000 1026.725000 0.630000 ;
      RECT 1017.415000 0.000000 1021.860000 0.630000 ;
      RECT 1012.545000 0.000000 1016.995000 0.630000 ;
      RECT 1007.680000 0.000000 1012.125000 0.630000 ;
      RECT 1002.810000 0.000000 1007.260000 0.630000 ;
      RECT 997.945000 0.000000 1002.390000 0.630000 ;
      RECT 993.080000 0.000000 997.525000 0.630000 ;
      RECT 988.210000 0.000000 992.660000 0.630000 ;
      RECT 983.345000 0.000000 987.790000 0.630000 ;
      RECT 978.475000 0.000000 982.925000 0.630000 ;
      RECT 973.610000 0.000000 978.055000 0.630000 ;
      RECT 968.745000 0.000000 973.190000 0.630000 ;
      RECT 963.875000 0.000000 968.325000 0.630000 ;
      RECT 959.010000 0.000000 963.455000 0.630000 ;
      RECT 954.140000 0.000000 958.590000 0.630000 ;
      RECT 949.275000 0.000000 953.720000 0.630000 ;
      RECT 944.410000 0.000000 948.855000 0.630000 ;
      RECT 939.540000 0.000000 943.990000 0.630000 ;
      RECT 934.675000 0.000000 939.120000 0.630000 ;
      RECT 929.805000 0.000000 934.255000 0.630000 ;
      RECT 924.940000 0.000000 929.385000 0.630000 ;
      RECT 920.075000 0.000000 924.520000 0.630000 ;
      RECT 915.205000 0.000000 919.655000 0.630000 ;
      RECT 910.340000 0.000000 914.785000 0.630000 ;
      RECT 905.470000 0.000000 909.920000 0.630000 ;
      RECT 900.605000 0.000000 905.050000 0.630000 ;
      RECT 895.740000 0.000000 900.185000 0.630000 ;
      RECT 890.870000 0.000000 895.320000 0.630000 ;
      RECT 886.005000 0.000000 890.450000 0.630000 ;
      RECT 881.135000 0.000000 885.585000 0.630000 ;
      RECT 876.270000 0.000000 880.715000 0.630000 ;
      RECT 871.405000 0.000000 875.850000 0.630000 ;
      RECT 866.535000 0.000000 870.985000 0.630000 ;
      RECT 861.670000 0.000000 866.115000 0.630000 ;
      RECT 856.800000 0.000000 861.250000 0.630000 ;
      RECT 851.935000 0.000000 856.380000 0.630000 ;
      RECT 847.070000 0.000000 851.515000 0.630000 ;
      RECT 842.200000 0.000000 846.650000 0.630000 ;
      RECT 837.335000 0.000000 841.780000 0.630000 ;
      RECT 832.465000 0.000000 836.915000 0.630000 ;
      RECT 827.600000 0.000000 832.045000 0.630000 ;
      RECT 822.735000 0.000000 827.180000 0.630000 ;
      RECT 817.865000 0.000000 822.315000 0.630000 ;
      RECT 813.000000 0.000000 817.445000 0.630000 ;
      RECT 808.130000 0.000000 812.580000 0.630000 ;
      RECT 803.265000 0.000000 807.710000 0.630000 ;
      RECT 798.400000 0.000000 802.845000 0.630000 ;
      RECT 793.530000 0.000000 797.980000 0.630000 ;
      RECT 788.665000 0.000000 793.110000 0.630000 ;
      RECT 783.795000 0.000000 788.245000 0.630000 ;
      RECT 778.930000 0.000000 783.375000 0.630000 ;
      RECT 774.065000 0.000000 778.510000 0.630000 ;
      RECT 769.195000 0.000000 773.645000 0.630000 ;
      RECT 764.330000 0.000000 768.775000 0.630000 ;
      RECT 759.460000 0.000000 763.910000 0.630000 ;
      RECT 754.595000 0.000000 759.040000 0.630000 ;
      RECT 749.730000 0.000000 754.175000 0.630000 ;
      RECT 744.860000 0.000000 749.310000 0.630000 ;
      RECT 739.995000 0.000000 744.440000 0.630000 ;
      RECT 735.125000 0.000000 739.575000 0.630000 ;
      RECT 730.260000 0.000000 734.705000 0.630000 ;
      RECT 725.395000 0.000000 729.840000 0.630000 ;
      RECT 720.525000 0.000000 724.975000 0.630000 ;
      RECT 715.660000 0.000000 720.105000 0.630000 ;
      RECT 710.790000 0.000000 715.240000 0.630000 ;
      RECT 705.925000 0.000000 710.370000 0.630000 ;
      RECT 701.060000 0.000000 705.505000 0.630000 ;
      RECT 696.190000 0.000000 700.640000 0.630000 ;
      RECT 691.325000 0.000000 695.770000 0.630000 ;
      RECT 686.455000 0.000000 690.905000 0.630000 ;
      RECT 681.590000 0.000000 686.035000 0.630000 ;
      RECT 676.725000 0.000000 681.170000 0.630000 ;
      RECT 671.855000 0.000000 676.305000 0.630000 ;
      RECT 666.990000 0.000000 671.435000 0.630000 ;
      RECT 662.120000 0.000000 666.570000 0.630000 ;
      RECT 657.255000 0.000000 661.700000 0.630000 ;
      RECT 652.390000 0.000000 656.835000 0.630000 ;
      RECT 647.520000 0.000000 651.970000 0.630000 ;
      RECT 642.655000 0.000000 647.100000 0.630000 ;
      RECT 637.785000 0.000000 642.235000 0.630000 ;
      RECT 632.920000 0.000000 637.365000 0.630000 ;
      RECT 628.055000 0.000000 632.500000 0.630000 ;
      RECT 623.185000 0.000000 627.635000 0.630000 ;
      RECT 618.320000 0.000000 622.765000 0.630000 ;
      RECT 613.450000 0.000000 617.900000 0.630000 ;
      RECT 608.585000 0.000000 613.030000 0.630000 ;
      RECT 603.720000 0.000000 608.165000 0.630000 ;
      RECT 598.850000 0.000000 603.300000 0.630000 ;
      RECT 593.985000 0.000000 598.430000 0.630000 ;
      RECT 589.115000 0.000000 593.565000 0.630000 ;
      RECT 584.250000 0.000000 588.695000 0.630000 ;
      RECT 579.385000 0.000000 583.830000 0.630000 ;
      RECT 574.515000 0.000000 578.965000 0.630000 ;
      RECT 569.650000 0.000000 574.095000 0.630000 ;
      RECT 564.780000 0.000000 569.230000 0.630000 ;
      RECT 559.915000 0.000000 564.360000 0.630000 ;
      RECT 555.050000 0.000000 559.495000 0.630000 ;
      RECT 550.180000 0.000000 554.630000 0.630000 ;
      RECT 545.315000 0.000000 549.760000 0.630000 ;
      RECT 540.445000 0.000000 544.895000 0.630000 ;
      RECT 535.580000 0.000000 540.025000 0.630000 ;
      RECT 530.715000 0.000000 535.160000 0.630000 ;
      RECT 525.845000 0.000000 530.295000 0.630000 ;
      RECT 520.980000 0.000000 525.425000 0.630000 ;
      RECT 516.110000 0.000000 520.560000 0.630000 ;
      RECT 511.245000 0.000000 515.690000 0.630000 ;
      RECT 506.380000 0.000000 510.825000 0.630000 ;
      RECT 501.510000 0.000000 505.960000 0.630000 ;
      RECT 496.645000 0.000000 501.090000 0.630000 ;
      RECT 491.775000 0.000000 496.225000 0.630000 ;
      RECT 486.910000 0.000000 491.355000 0.630000 ;
      RECT 482.045000 0.000000 486.490000 0.630000 ;
      RECT 477.175000 0.000000 481.625000 0.630000 ;
      RECT 472.310000 0.000000 476.755000 0.630000 ;
      RECT 467.440000 0.000000 471.890000 0.630000 ;
      RECT 462.575000 0.000000 467.020000 0.630000 ;
      RECT 457.710000 0.000000 462.155000 0.630000 ;
      RECT 452.840000 0.000000 457.290000 0.630000 ;
      RECT 447.975000 0.000000 452.420000 0.630000 ;
      RECT 443.105000 0.000000 447.555000 0.630000 ;
      RECT 438.240000 0.000000 442.685000 0.630000 ;
      RECT 433.375000 0.000000 437.820000 0.630000 ;
      RECT 428.505000 0.000000 432.955000 0.630000 ;
      RECT 423.640000 0.000000 428.085000 0.630000 ;
      RECT 418.770000 0.000000 423.220000 0.630000 ;
      RECT 413.905000 0.000000 418.350000 0.630000 ;
      RECT 409.040000 0.000000 413.485000 0.630000 ;
      RECT 404.170000 0.000000 408.620000 0.630000 ;
      RECT 399.305000 0.000000 403.750000 0.630000 ;
      RECT 394.435000 0.000000 398.885000 0.630000 ;
      RECT 389.570000 0.000000 394.015000 0.630000 ;
      RECT 384.705000 0.000000 389.150000 0.630000 ;
      RECT 379.835000 0.000000 384.285000 0.630000 ;
      RECT 374.970000 0.000000 379.415000 0.630000 ;
      RECT 370.100000 0.000000 374.550000 0.630000 ;
      RECT 365.235000 0.000000 369.680000 0.630000 ;
      RECT 360.370000 0.000000 364.815000 0.630000 ;
      RECT 355.500000 0.000000 359.950000 0.630000 ;
      RECT 350.635000 0.000000 355.080000 0.630000 ;
      RECT 345.765000 0.000000 350.215000 0.630000 ;
      RECT 340.900000 0.000000 345.345000 0.630000 ;
      RECT 336.035000 0.000000 340.480000 0.630000 ;
      RECT 331.165000 0.000000 335.615000 0.630000 ;
      RECT 326.300000 0.000000 330.745000 0.630000 ;
      RECT 321.430000 0.000000 325.880000 0.630000 ;
      RECT 316.565000 0.000000 321.010000 0.630000 ;
      RECT 311.700000 0.000000 316.145000 0.630000 ;
      RECT 306.830000 0.000000 311.280000 0.630000 ;
      RECT 301.965000 0.000000 306.410000 0.630000 ;
      RECT 297.095000 0.000000 301.545000 0.630000 ;
      RECT 292.230000 0.000000 296.675000 0.630000 ;
      RECT 287.365000 0.000000 291.810000 0.630000 ;
      RECT 282.495000 0.000000 286.945000 0.630000 ;
      RECT 277.630000 0.000000 282.075000 0.630000 ;
      RECT 272.760000 0.000000 277.210000 0.630000 ;
      RECT 267.895000 0.000000 272.340000 0.630000 ;
      RECT 263.030000 0.000000 267.475000 0.630000 ;
      RECT 258.160000 0.000000 262.610000 0.630000 ;
      RECT 253.295000 0.000000 257.740000 0.630000 ;
      RECT 248.425000 0.000000 252.875000 0.630000 ;
      RECT 243.560000 0.000000 248.005000 0.630000 ;
      RECT 238.695000 0.000000 243.140000 0.630000 ;
      RECT 233.825000 0.000000 238.275000 0.630000 ;
      RECT 228.960000 0.000000 233.405000 0.630000 ;
      RECT 224.090000 0.000000 228.540000 0.630000 ;
      RECT 219.225000 0.000000 223.670000 0.630000 ;
      RECT 214.360000 0.000000 218.805000 0.630000 ;
      RECT 209.490000 0.000000 213.940000 0.630000 ;
      RECT 204.625000 0.000000 209.070000 0.630000 ;
      RECT 199.755000 0.000000 204.205000 0.630000 ;
      RECT 194.890000 0.000000 199.335000 0.630000 ;
      RECT 190.025000 0.000000 194.470000 0.630000 ;
      RECT 185.155000 0.000000 189.605000 0.630000 ;
      RECT 180.290000 0.000000 184.735000 0.630000 ;
      RECT 175.420000 0.000000 179.870000 0.630000 ;
      RECT 170.555000 0.000000 175.000000 0.630000 ;
      RECT 165.690000 0.000000 170.135000 0.630000 ;
      RECT 160.820000 0.000000 165.270000 0.630000 ;
      RECT 155.955000 0.000000 160.400000 0.630000 ;
      RECT 151.085000 0.000000 155.535000 0.630000 ;
      RECT 146.220000 0.000000 150.665000 0.630000 ;
      RECT 141.355000 0.000000 145.800000 0.630000 ;
      RECT 136.485000 0.000000 140.935000 0.630000 ;
      RECT 131.620000 0.000000 136.065000 0.630000 ;
      RECT 126.750000 0.000000 131.200000 0.630000 ;
      RECT 121.885000 0.000000 126.330000 0.630000 ;
      RECT 117.020000 0.000000 121.465000 0.630000 ;
      RECT 112.150000 0.000000 116.600000 0.630000 ;
      RECT 107.285000 0.000000 111.730000 0.630000 ;
      RECT 102.415000 0.000000 106.865000 0.630000 ;
      RECT 97.550000 0.000000 101.995000 0.630000 ;
      RECT 92.685000 0.000000 97.130000 0.630000 ;
      RECT 87.815000 0.000000 92.265000 0.630000 ;
      RECT 82.950000 0.000000 87.395000 0.630000 ;
      RECT 78.080000 0.000000 82.530000 0.630000 ;
      RECT 73.215000 0.000000 77.660000 0.630000 ;
      RECT 68.350000 0.000000 72.795000 0.630000 ;
      RECT 63.480000 0.000000 67.930000 0.630000 ;
      RECT 58.615000 0.000000 63.060000 0.630000 ;
      RECT 53.745000 0.000000 58.195000 0.630000 ;
      RECT 48.880000 0.000000 53.325000 0.630000 ;
      RECT 44.015000 0.000000 48.460000 0.630000 ;
      RECT 39.145000 0.000000 43.595000 0.630000 ;
      RECT 34.280000 0.000000 38.725000 0.630000 ;
      RECT 29.410000 0.000000 33.860000 0.630000 ;
      RECT 24.545000 0.000000 28.990000 0.630000 ;
      RECT 19.680000 0.000000 24.125000 0.630000 ;
      RECT 14.810000 0.000000 19.260000 0.630000 ;
      RECT 9.945000 0.000000 14.390000 0.630000 ;
      RECT 5.075000 0.000000 9.525000 0.630000 ;
      RECT 0.000000 0.000000 4.655000 0.630000 ;
    LAYER met3 ;
      RECT 0.000000 2599.930000 2399.820000 2599.980000 ;
      RECT 0.000000 2599.030000 2398.720000 2599.930000 ;
      RECT 0.000000 2598.710000 2399.820000 2599.030000 ;
      RECT 1.100000 2597.810000 2399.820000 2598.710000 ;
      RECT 0.000000 2551.360000 2399.820000 2597.810000 ;
      RECT 1.100000 2550.460000 2399.820000 2551.360000 ;
      RECT 0.000000 2550.400000 2399.820000 2550.460000 ;
      RECT 0.000000 2549.500000 2398.720000 2550.400000 ;
      RECT 0.000000 2502.305000 2399.820000 2549.500000 ;
      RECT 1.100000 2501.405000 2399.820000 2502.305000 ;
      RECT 0.000000 2500.400000 2399.820000 2501.405000 ;
      RECT 0.000000 2499.500000 2398.720000 2500.400000 ;
      RECT 0.000000 2453.250000 2399.820000 2499.500000 ;
      RECT 1.100000 2452.350000 2399.820000 2453.250000 ;
      RECT 0.000000 2450.400000 2399.820000 2452.350000 ;
      RECT 0.000000 2449.500000 2398.720000 2450.400000 ;
      RECT 0.000000 2404.195000 2399.820000 2449.500000 ;
      RECT 1.100000 2403.295000 2399.820000 2404.195000 ;
      RECT 0.000000 2400.400000 2399.820000 2403.295000 ;
      RECT 0.000000 2399.500000 2398.720000 2400.400000 ;
      RECT 0.000000 2355.140000 2399.820000 2399.500000 ;
      RECT 1.100000 2354.240000 2399.820000 2355.140000 ;
      RECT 0.000000 2350.405000 2399.820000 2354.240000 ;
      RECT 0.000000 2349.505000 2398.720000 2350.405000 ;
      RECT 0.000000 2306.080000 2399.820000 2349.505000 ;
      RECT 1.100000 2305.180000 2399.820000 2306.080000 ;
      RECT 0.000000 2300.405000 2399.820000 2305.180000 ;
      RECT 0.000000 2299.505000 2398.720000 2300.405000 ;
      RECT 0.000000 2257.025000 2399.820000 2299.505000 ;
      RECT 1.100000 2256.125000 2399.820000 2257.025000 ;
      RECT 0.000000 2250.405000 2399.820000 2256.125000 ;
      RECT 0.000000 2249.505000 2398.720000 2250.405000 ;
      RECT 0.000000 2207.970000 2399.820000 2249.505000 ;
      RECT 1.100000 2207.070000 2399.820000 2207.970000 ;
      RECT 0.000000 2200.405000 2399.820000 2207.070000 ;
      RECT 0.000000 2199.505000 2398.720000 2200.405000 ;
      RECT 0.000000 2158.915000 2399.820000 2199.505000 ;
      RECT 1.100000 2158.015000 2399.820000 2158.915000 ;
      RECT 0.000000 2150.405000 2399.820000 2158.015000 ;
      RECT 0.000000 2149.505000 2398.720000 2150.405000 ;
      RECT 0.000000 2109.860000 2399.820000 2149.505000 ;
      RECT 1.100000 2108.960000 2399.820000 2109.860000 ;
      RECT 0.000000 2100.410000 2399.820000 2108.960000 ;
      RECT 0.000000 2099.510000 2398.720000 2100.410000 ;
      RECT 0.000000 2060.800000 2399.820000 2099.510000 ;
      RECT 1.100000 2059.900000 2399.820000 2060.800000 ;
      RECT 0.000000 2050.410000 2399.820000 2059.900000 ;
      RECT 0.000000 2049.510000 2398.720000 2050.410000 ;
      RECT 0.000000 2011.745000 2399.820000 2049.510000 ;
      RECT 1.100000 2010.845000 2399.820000 2011.745000 ;
      RECT 0.000000 2000.410000 2399.820000 2010.845000 ;
      RECT 0.000000 1999.510000 2398.720000 2000.410000 ;
      RECT 0.000000 1962.690000 2399.820000 1999.510000 ;
      RECT 1.100000 1961.790000 2399.820000 1962.690000 ;
      RECT 0.000000 1950.410000 2399.820000 1961.790000 ;
      RECT 0.000000 1949.510000 2398.720000 1950.410000 ;
      RECT 0.000000 1913.635000 2399.820000 1949.510000 ;
      RECT 1.100000 1912.735000 2399.820000 1913.635000 ;
      RECT 0.000000 1900.410000 2399.820000 1912.735000 ;
      RECT 0.000000 1899.510000 2398.720000 1900.410000 ;
      RECT 0.000000 1864.580000 2399.820000 1899.510000 ;
      RECT 1.100000 1863.680000 2399.820000 1864.580000 ;
      RECT 0.000000 1850.415000 2399.820000 1863.680000 ;
      RECT 0.000000 1849.515000 2398.720000 1850.415000 ;
      RECT 0.000000 1815.520000 2399.820000 1849.515000 ;
      RECT 1.100000 1814.620000 2399.820000 1815.520000 ;
      RECT 0.000000 1800.415000 2399.820000 1814.620000 ;
      RECT 0.000000 1799.515000 2398.720000 1800.415000 ;
      RECT 0.000000 1766.465000 2399.820000 1799.515000 ;
      RECT 1.100000 1765.565000 2399.820000 1766.465000 ;
      RECT 0.000000 1750.415000 2399.820000 1765.565000 ;
      RECT 0.000000 1749.515000 2398.720000 1750.415000 ;
      RECT 0.000000 1717.410000 2399.820000 1749.515000 ;
      RECT 1.100000 1716.510000 2399.820000 1717.410000 ;
      RECT 0.000000 1700.415000 2399.820000 1716.510000 ;
      RECT 0.000000 1699.515000 2398.720000 1700.415000 ;
      RECT 0.000000 1668.355000 2399.820000 1699.515000 ;
      RECT 1.100000 1667.455000 2399.820000 1668.355000 ;
      RECT 0.000000 1650.415000 2399.820000 1667.455000 ;
      RECT 0.000000 1649.515000 2398.720000 1650.415000 ;
      RECT 0.000000 1619.300000 2399.820000 1649.515000 ;
      RECT 1.100000 1618.400000 2399.820000 1619.300000 ;
      RECT 0.000000 1600.420000 2399.820000 1618.400000 ;
      RECT 0.000000 1599.520000 2398.720000 1600.420000 ;
      RECT 0.000000 1570.240000 2399.820000 1599.520000 ;
      RECT 1.100000 1569.340000 2399.820000 1570.240000 ;
      RECT 0.000000 1550.420000 2399.820000 1569.340000 ;
      RECT 0.000000 1549.520000 2398.720000 1550.420000 ;
      RECT 0.000000 1521.185000 2399.820000 1549.520000 ;
      RECT 1.100000 1520.285000 2399.820000 1521.185000 ;
      RECT 0.000000 1500.420000 2399.820000 1520.285000 ;
      RECT 0.000000 1499.520000 2398.720000 1500.420000 ;
      RECT 0.000000 1472.130000 2399.820000 1499.520000 ;
      RECT 1.100000 1471.230000 2399.820000 1472.130000 ;
      RECT 0.000000 1450.420000 2399.820000 1471.230000 ;
      RECT 0.000000 1449.520000 2398.720000 1450.420000 ;
      RECT 0.000000 1423.075000 2399.820000 1449.520000 ;
      RECT 1.100000 1422.175000 2399.820000 1423.075000 ;
      RECT 0.000000 1400.420000 2399.820000 1422.175000 ;
      RECT 0.000000 1399.520000 2398.720000 1400.420000 ;
      RECT 0.000000 1374.020000 2399.820000 1399.520000 ;
      RECT 1.100000 1373.120000 2399.820000 1374.020000 ;
      RECT 0.000000 1350.425000 2399.820000 1373.120000 ;
      RECT 0.000000 1349.525000 2398.720000 1350.425000 ;
      RECT 0.000000 1324.960000 2399.820000 1349.525000 ;
      RECT 1.100000 1324.060000 2399.820000 1324.960000 ;
      RECT 0.000000 1300.425000 2399.820000 1324.060000 ;
      RECT 0.000000 1299.525000 2398.720000 1300.425000 ;
      RECT 0.000000 1275.905000 2399.820000 1299.525000 ;
      RECT 1.100000 1275.005000 2399.820000 1275.905000 ;
      RECT 0.000000 1250.425000 2399.820000 1275.005000 ;
      RECT 0.000000 1249.525000 2398.720000 1250.425000 ;
      RECT 0.000000 1226.850000 2399.820000 1249.525000 ;
      RECT 1.100000 1225.950000 2399.820000 1226.850000 ;
      RECT 0.000000 1200.425000 2399.820000 1225.950000 ;
      RECT 0.000000 1199.525000 2398.720000 1200.425000 ;
      RECT 0.000000 1177.795000 2399.820000 1199.525000 ;
      RECT 1.100000 1176.895000 2399.820000 1177.795000 ;
      RECT 0.000000 1150.425000 2399.820000 1176.895000 ;
      RECT 0.000000 1149.525000 2398.720000 1150.425000 ;
      RECT 0.000000 1128.740000 2399.820000 1149.525000 ;
      RECT 1.100000 1127.840000 2399.820000 1128.740000 ;
      RECT 0.000000 1100.430000 2399.820000 1127.840000 ;
      RECT 0.000000 1099.530000 2398.720000 1100.430000 ;
      RECT 0.000000 1079.680000 2399.820000 1099.530000 ;
      RECT 1.100000 1078.780000 2399.820000 1079.680000 ;
      RECT 0.000000 1050.430000 2399.820000 1078.780000 ;
      RECT 0.000000 1049.530000 2398.720000 1050.430000 ;
      RECT 0.000000 1030.625000 2399.820000 1049.530000 ;
      RECT 1.100000 1029.725000 2399.820000 1030.625000 ;
      RECT 0.000000 1000.430000 2399.820000 1029.725000 ;
      RECT 0.000000 999.530000 2398.720000 1000.430000 ;
      RECT 0.000000 981.570000 2399.820000 999.530000 ;
      RECT 1.100000 980.670000 2399.820000 981.570000 ;
      RECT 0.000000 950.430000 2399.820000 980.670000 ;
      RECT 0.000000 949.530000 2398.720000 950.430000 ;
      RECT 0.000000 932.515000 2399.820000 949.530000 ;
      RECT 1.100000 931.615000 2399.820000 932.515000 ;
      RECT 0.000000 900.430000 2399.820000 931.615000 ;
      RECT 0.000000 899.530000 2398.720000 900.430000 ;
      RECT 0.000000 883.460000 2399.820000 899.530000 ;
      RECT 1.100000 882.560000 2399.820000 883.460000 ;
      RECT 0.000000 850.435000 2399.820000 882.560000 ;
      RECT 0.000000 849.535000 2398.720000 850.435000 ;
      RECT 0.000000 834.400000 2399.820000 849.535000 ;
      RECT 1.100000 833.500000 2399.820000 834.400000 ;
      RECT 0.000000 800.435000 2399.820000 833.500000 ;
      RECT 0.000000 799.535000 2398.720000 800.435000 ;
      RECT 0.000000 785.345000 2399.820000 799.535000 ;
      RECT 1.100000 784.445000 2399.820000 785.345000 ;
      RECT 0.000000 750.435000 2399.820000 784.445000 ;
      RECT 0.000000 749.535000 2398.720000 750.435000 ;
      RECT 0.000000 736.290000 2399.820000 749.535000 ;
      RECT 1.100000 735.390000 2399.820000 736.290000 ;
      RECT 0.000000 700.435000 2399.820000 735.390000 ;
      RECT 0.000000 699.535000 2398.720000 700.435000 ;
      RECT 0.000000 687.235000 2399.820000 699.535000 ;
      RECT 1.100000 686.335000 2399.820000 687.235000 ;
      RECT 0.000000 650.435000 2399.820000 686.335000 ;
      RECT 0.000000 649.535000 2398.720000 650.435000 ;
      RECT 0.000000 638.180000 2399.820000 649.535000 ;
      RECT 1.100000 637.280000 2399.820000 638.180000 ;
      RECT 0.000000 600.440000 2399.820000 637.280000 ;
      RECT 0.000000 599.540000 2398.720000 600.440000 ;
      RECT 0.000000 589.120000 2399.820000 599.540000 ;
      RECT 1.100000 588.220000 2399.820000 589.120000 ;
      RECT 0.000000 550.440000 2399.820000 588.220000 ;
      RECT 0.000000 549.540000 2398.720000 550.440000 ;
      RECT 0.000000 540.065000 2399.820000 549.540000 ;
      RECT 1.100000 539.165000 2399.820000 540.065000 ;
      RECT 0.000000 500.440000 2399.820000 539.165000 ;
      RECT 0.000000 499.540000 2398.720000 500.440000 ;
      RECT 0.000000 491.010000 2399.820000 499.540000 ;
      RECT 1.100000 490.110000 2399.820000 491.010000 ;
      RECT 0.000000 450.440000 2399.820000 490.110000 ;
      RECT 0.000000 449.540000 2398.720000 450.440000 ;
      RECT 0.000000 441.955000 2399.820000 449.540000 ;
      RECT 1.100000 441.055000 2399.820000 441.955000 ;
      RECT 0.000000 400.440000 2399.820000 441.055000 ;
      RECT 0.000000 399.540000 2398.720000 400.440000 ;
      RECT 0.000000 392.900000 2399.820000 399.540000 ;
      RECT 1.100000 392.000000 2399.820000 392.900000 ;
      RECT 0.000000 350.445000 2399.820000 392.000000 ;
      RECT 0.000000 349.545000 2398.720000 350.445000 ;
      RECT 0.000000 343.840000 2399.820000 349.545000 ;
      RECT 1.100000 342.940000 2399.820000 343.840000 ;
      RECT 0.000000 300.445000 2399.820000 342.940000 ;
      RECT 0.000000 299.545000 2398.720000 300.445000 ;
      RECT 0.000000 294.785000 2399.820000 299.545000 ;
      RECT 1.100000 293.885000 2399.820000 294.785000 ;
      RECT 0.000000 250.445000 2399.820000 293.885000 ;
      RECT 0.000000 249.545000 2398.720000 250.445000 ;
      RECT 0.000000 245.730000 2399.820000 249.545000 ;
      RECT 1.100000 244.830000 2399.820000 245.730000 ;
      RECT 0.000000 200.445000 2399.820000 244.830000 ;
      RECT 0.000000 199.545000 2398.720000 200.445000 ;
      RECT 0.000000 196.675000 2399.820000 199.545000 ;
      RECT 1.100000 195.775000 2399.820000 196.675000 ;
      RECT 0.000000 150.445000 2399.820000 195.775000 ;
      RECT 0.000000 149.545000 2398.720000 150.445000 ;
      RECT 0.000000 147.620000 2399.820000 149.545000 ;
      RECT 1.100000 146.720000 2399.820000 147.620000 ;
      RECT 0.000000 100.450000 2399.820000 146.720000 ;
      RECT 0.000000 99.550000 2398.720000 100.450000 ;
      RECT 0.000000 98.560000 2399.820000 99.550000 ;
      RECT 1.100000 97.660000 2399.820000 98.560000 ;
      RECT 0.000000 50.450000 2399.820000 97.660000 ;
      RECT 0.000000 49.550000 2398.720000 50.450000 ;
      RECT 0.000000 49.505000 2399.820000 49.550000 ;
      RECT 1.100000 48.605000 2399.820000 49.505000 ;
      RECT 0.000000 3.770000 2399.820000 48.605000 ;
      RECT 0.000000 2.870000 2398.720000 3.770000 ;
      RECT 0.000000 1.100000 2399.820000 2.870000 ;
      RECT 2.060000 0.000000 2399.820000 1.100000 ;
      RECT 0.000000 0.000000 1.160000 1.100000 ;
    LAYER met4 ;
      RECT 0.000000 2595.920000 2399.820000 2599.980000 ;
      RECT 5.020000 2592.320000 2394.800000 2595.920000 ;
      RECT 8.620000 2592.300000 2394.800000 2592.320000 ;
      RECT 2393.600000 5.960000 2394.800000 2592.300000 ;
      RECT 8.620000 5.960000 2391.260000 2592.300000 ;
      RECT 5.020000 5.960000 6.220000 2592.320000 ;
      RECT 2397.200000 2.360000 2399.820000 2595.920000 ;
      RECT 5.020000 2.360000 2394.800000 5.960000 ;
      RECT 0.000000 2.360000 2.620000 2595.920000 ;
      RECT 0.000000 0.000000 2399.820000 2.360000 ;
    LAYER met5 ;
      RECT 0.000000 0.000000 2399.820000 2599.980000 ;
  END
END azadi_soc_top_caravel

END LIBRARY
